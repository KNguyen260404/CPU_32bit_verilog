* NGSPICE file created from CPU_core.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_2 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

.subckt CPU_core VGND VPWR clk debug_reg1[0] debug_reg1[10] debug_reg1[11] debug_reg1[12]
+ debug_reg1[13] debug_reg1[14] debug_reg1[15] debug_reg1[16] debug_reg1[17] debug_reg1[18]
+ debug_reg1[19] debug_reg1[1] debug_reg1[20] debug_reg1[21] debug_reg1[22] debug_reg1[23]
+ debug_reg1[24] debug_reg1[25] debug_reg1[26] debug_reg1[27] debug_reg1[28] debug_reg1[29]
+ debug_reg1[2] debug_reg1[30] debug_reg1[31] debug_reg1[3] debug_reg1[4] debug_reg1[5]
+ debug_reg1[6] debug_reg1[7] debug_reg1[8] debug_reg1[9] debug_reg2[0] debug_reg2[10]
+ debug_reg2[11] debug_reg2[12] debug_reg2[13] debug_reg2[14] debug_reg2[15] debug_reg2[16]
+ debug_reg2[17] debug_reg2[18] debug_reg2[19] debug_reg2[1] debug_reg2[20] debug_reg2[21]
+ debug_reg2[22] debug_reg2[23] debug_reg2[24] debug_reg2[25] debug_reg2[26] debug_reg2[27]
+ debug_reg2[28] debug_reg2[29] debug_reg2[2] debug_reg2[30] debug_reg2[31] debug_reg2[3]
+ debug_reg2[4] debug_reg2[5] debug_reg2[6] debug_reg2[7] debug_reg2[8] debug_reg2[9]
+ debug_reg3[0] debug_reg3[10] debug_reg3[11] debug_reg3[12] debug_reg3[13] debug_reg3[14]
+ debug_reg3[15] debug_reg3[16] debug_reg3[17] debug_reg3[18] debug_reg3[19] debug_reg3[1]
+ debug_reg3[20] debug_reg3[21] debug_reg3[22] debug_reg3[23] debug_reg3[24] debug_reg3[25]
+ debug_reg3[26] debug_reg3[27] debug_reg3[28] debug_reg3[29] debug_reg3[2] debug_reg3[30]
+ debug_reg3[31] debug_reg3[3] debug_reg3[4] debug_reg3[5] debug_reg3[6] debug_reg3[7]
+ debug_reg3[8] debug_reg3[9] instruction_debug[0] instruction_debug[10] instruction_debug[11]
+ instruction_debug[12] instruction_debug[13] instruction_debug[14] instruction_debug[15]
+ instruction_debug[16] instruction_debug[17] instruction_debug[18] instruction_debug[19]
+ instruction_debug[1] instruction_debug[20] instruction_debug[21] instruction_debug[22]
+ instruction_debug[23] instruction_debug[27] instruction_debug[2] instruction_debug[30]
+ instruction_debug[31] instruction_debug[3] instruction_debug[4] instruction_debug[5]
+ instruction_debug[6] instruction_debug[7] instruction_debug[8] instruction_debug[9]
+ pc_current[0] pc_current[10] pc_current[11] pc_current[12] pc_current[13] pc_current[14]
+ pc_current[15] pc_current[16] pc_current[17] pc_current[18] pc_current[19] pc_current[1]
+ pc_current[20] pc_current[21] pc_current[22] pc_current[23] pc_current[24] pc_current[25]
+ pc_current[26] pc_current[27] pc_current[28] pc_current[29] pc_current[2] pc_current[30]
+ pc_current[31] pc_current[3] pc_current[4] pc_current[5] pc_current[6] pc_current[7]
+ pc_current[8] pc_current[9] pipeline_state[0] pipeline_state[1] pipeline_state[2]
+ pipeline_state[3] reset instruction_debug[26] instruction_debug[25] instruction_debug[24]
+ instruction_debug[29] instruction_debug[28]
XFILLER_0_89_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold340 net17 VGND VGND VPWR VPWR net535 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1270_ _0307_ _0309_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_17_Left_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0985_ _0623_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XCPU_core_149 VGND VGND VPWR VPWR CPU_core_149/HI instruction_debug[12] sky130_fd_sc_hd__conb_1
XFILLER_0_42_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1606_ net300 _0512_ _0514_ net483 VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_26_Left_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1537_ net366 _0503_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__and2_1
X_1468_ net512 _0478_ _0480_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__o21a_1
X_1399_ _0519_ net490 VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_2_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold170 net4 VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 net66 VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 dmem.address\[16\] VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1322_ _0837_ _0375_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__nand2_1
X_1253_ _0310_ _0311_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1184_ dmem.address\[18\] _0809_ _0611_ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_86_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0968_ _0603_ _0605_ _0607_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_113_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0899_ net395 VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1940_ clknet_leaf_3_clk _0256_ VGND VGND VPWR VPWR id_ex_rs1_data\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1871_ clknet_leaf_2_clk net263 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_87 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1305_ _0329_ _0334_ _0342_ _0357_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__a211o_1
X_1236_ _0773_ _0832_ _0838_ _0293_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__o31a_1
XFILLER_0_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1167_ _0594_ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1098_ _0711_ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1021_ _0648_ _0650_ _0656_ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_37_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1923_ clknet_leaf_19_clk _0239_ VGND VGND VPWR VPWR id_alu_src\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1854_ clknet_leaf_8_clk _0170_ VGND VGND VPWR VPWR id_ex_rs2_data\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1785_ clknet_leaf_12_clk net513 VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_762 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1219_ net335 _0556_ _0279_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold41 net72 VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 _0227_ VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 _0122_ VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 _0190_ VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 net30 VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold85 register_file.write_data\[26\] VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 _0175_ VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1570_ net290 _0506_ _0508_ net55 VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1004_ _0628_ _0640_ _0641_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1906_ clknet_leaf_1_clk net215 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_114_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1837_ clknet_leaf_2_clk _0153_ VGND VGND VPWR VPWR id_ex_rs2_data\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1768_ clknet_leaf_14_clk _0084_ VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1699_ clknet_leaf_3_clk _0016_ VGND VGND VPWR VPWR register_file.write_data\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_99_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput42 net42 VGND VGND VPWR VPWR debug_reg2[18] sky130_fd_sc_hd__buf_8
Xoutput31 net31 VGND VGND VPWR VPWR debug_reg1[8] sky130_fd_sc_hd__buf_8
Xoutput7 net7 VGND VGND VPWR VPWR debug_reg1[15] sky130_fd_sc_hd__buf_12
XFILLER_0_31_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput20 net20 VGND VGND VPWR VPWR debug_reg1[27] sky130_fd_sc_hd__buf_8
XFILLER_0_101_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput75 net75 VGND VGND VPWR VPWR debug_reg3[19] sky130_fd_sc_hd__buf_8
Xoutput53 net53 VGND VGND VPWR VPWR debug_reg2[28] sky130_fd_sc_hd__buf_8
Xoutput64 net64 VGND VGND VPWR VPWR debug_reg2[9] sky130_fd_sc_hd__buf_8
Xoutput86 net86 VGND VGND VPWR VPWR debug_reg3[29] sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_8_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput97 net97 VGND VGND VPWR VPWR instruction_debug[15] sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_47_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1622_ net208 _0515_ _0516_ net6 VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1553_ net316 _0504_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1484_ _0607_ _0490_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_99_Left_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold341 register_file.write_data\[29\] VGND VGND VPWR VPWR net536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold330 net129 VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0984_ _0616_ _0617_ _0621_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__nor3_1
XFILLER_0_42_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1605_ _0513_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1536_ net488 _0503_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1467_ net512 _0478_ _0452_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_2_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1398_ _0441_ _0628_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_118_Right_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold160 net21 VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold171 net61 VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 net67 VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 _0017_ VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1321_ net200 _0374_ _0835_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__mux2_1
X_1252_ _0307_ _0309_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__or2_1
X_1183_ register_file.write_data\[18\] id_ex_rs2_data\[18\] _0609_ VGND VGND VPWR
+ VPWR _0809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0967_ _0521_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__buf_1
XFILLER_0_42_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0898_ _0526_ _0541_ id_ex_rs2_data\[0\] VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__o21a_1
XFILLER_0_112_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1519_ net224 _0500_ _0501_ net248 VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Left_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1870_ clknet_leaf_2_clk net275 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_54_Left_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1304_ _0358_ _0359_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_63_Left_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1235_ _0773_ _0832_ _0294_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_126_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1166_ _0765_ _0752_ _0720_ _0646_ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_126_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1097_ _0689_ _0693_ _0712_ VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1020_ _0632_ _0634_ _0652_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_37_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1922_ clknet_leaf_18_clk _0238_ VGND VGND VPWR VPWR id_reg_write sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1853_ clknet_leaf_8_clk _0169_ VGND VGND VPWR VPWR id_ex_rs2_data\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_54 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1784_ clknet_leaf_12_clk net450 VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_71_Left_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1218_ id_ex_rs1_data\[20\] _0558_ _0841_ _0532_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1149_ _0773_ _0776_ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_80_Left_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold20 _0222_ VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 register_file.write_data\[21\] VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 net79 VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 _0125_ VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 _0247_ VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold86 _0135_ VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 net34 VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 register_file.write_data\[3\] VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_119_Left_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_128_Left_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1003_ _0637_ _0639_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1905_ clknet_leaf_1_clk net207 VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dfxtp_2
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1836_ clknet_leaf_2_clk _0152_ VGND VGND VPWR VPWR id_ex_rs2_data\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1767_ clknet_leaf_14_clk _0083_ VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1698_ clknet_leaf_3_clk _0015_ VGND VGND VPWR VPWR register_file.write_data\[14\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_123_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput43 net43 VGND VGND VPWR VPWR debug_reg2[19] sky130_fd_sc_hd__buf_8
Xoutput32 net32 VGND VGND VPWR VPWR debug_reg1[9] sky130_fd_sc_hd__buf_8
XFILLER_0_31_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput8 net8 VGND VGND VPWR VPWR debug_reg1[16] sky130_fd_sc_hd__buf_12
Xoutput10 net10 VGND VGND VPWR VPWR debug_reg1[18] sky130_fd_sc_hd__buf_12
Xoutput21 net21 VGND VGND VPWR VPWR debug_reg1[28] sky130_fd_sc_hd__buf_8
XFILLER_0_101_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput76 net76 VGND VGND VPWR VPWR debug_reg3[1] sky130_fd_sc_hd__buf_8
Xoutput65 net65 VGND VGND VPWR VPWR debug_reg3[0] sky130_fd_sc_hd__buf_8
Xoutput54 net54 VGND VGND VPWR VPWR debug_reg2[29] sky130_fd_sc_hd__buf_8
Xoutput87 net87 VGND VGND VPWR VPWR debug_reg3[2] sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_8_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput98 net98 VGND VGND VPWR VPWR instruction_debug[20] sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_47_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1621_ net220 _0515_ _0516_ net5 VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1552_ net320 _0504_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1483_ net484 net479 _0487_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1819_ clknet_leaf_9_clk net281 VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dfxtp_1
Xhold320 _0092_ VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold342 net63 VGND VGND VPWR VPWR net537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 id_ex_immediate\[1\] VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0983_ _0616_ _0617_ _0621_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1604_ _0521_ net309 VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__nor2_4
XFILLER_0_10_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1535_ net389 _0503_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1466_ net449 _0477_ _0479_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__o21a_1
X_1397_ net337 VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__buf_2
XFILLER_0_97_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold161 _0268_ VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold150 net22 VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold183 register_file.write_data\[31\] VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 _0147_ VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 net59 VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1320_ register_file.write_data\[27\] id_ex_rs2_data\[27\] _0833_ VGND VGND VPWR
+ VPWR _0374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_775 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1251_ _0307_ _0309_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__nand2_1
X_1182_ _0807_ _0808_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0966_ _0603_ _0605_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0897_ forwarding_unit.rd_wb\[0\] forwarding_unit.rs2_ex\[3\] forwarding_unit.rs2_ex\[0\]
+ forwarding_unit.rs2_ex\[1\] VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__or4b_2
XFILLER_0_42_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1518_ net226 _0500_ _0501_ net286 VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1449_ _0452_ _0468_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_100_Left_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1303_ _0345_ _0344_ _0357_ _0607_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__a31o_1
X_1234_ _0838_ _0293_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_88_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1165_ _0628_ _0791_ _0792_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1096_ _0694_ _0698_ _0711_ _0712_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__nand4_1
XFILLER_0_87_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0949_ _0573_ _0575_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__and2b_1
XFILLER_0_43_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1921_ clknet_leaf_19_clk _0237_ VGND VGND VPWR VPWR forwarding_unit.reg_write_mem
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1852_ clknet_leaf_8_clk net348 VGND VGND VPWR VPWR id_ex_rs2_data\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1783_ clknet_leaf_12_clk net428 VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1217_ register_file.write_data\[20\] _0528_ VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__or2_1
X_1148_ _0594_ _0774_ _0775_ _0613_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1079_ _0707_ _0708_ _0710_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__or3_1
XFILLER_0_75_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold32 _0226_ VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 _0220_ VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 register_file.write_data\[18\] VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 _0131_ VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 net71 VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 net29 VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold87 register_file.write_data\[24\] VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 _0183_ VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 _0176_ VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_26 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1002_ _0637_ _0639_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1904_ clknet_leaf_1_clk net205 VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_127_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1835_ clknet_leaf_2_clk _0151_ VGND VGND VPWR VPWR id_ex_rs2_data\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_96_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1766_ clknet_leaf_15_clk net403 VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1697_ clknet_leaf_3_clk _0014_ VGND VGND VPWR VPWR register_file.write_data\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput9 net9 VGND VGND VPWR VPWR debug_reg1[17] sky130_fd_sc_hd__buf_12
Xoutput11 net11 VGND VGND VPWR VPWR debug_reg1[19] sky130_fd_sc_hd__buf_12
Xoutput22 net22 VGND VGND VPWR VPWR debug_reg1[29] sky130_fd_sc_hd__buf_8
Xoutput33 net33 VGND VGND VPWR VPWR debug_reg2[0] sky130_fd_sc_hd__buf_12
Xoutput66 net66 VGND VGND VPWR VPWR debug_reg3[10] sky130_fd_sc_hd__buf_8
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput44 net44 VGND VGND VPWR VPWR debug_reg2[1] sky130_fd_sc_hd__buf_12
Xoutput55 net55 VGND VGND VPWR VPWR debug_reg2[2] sky130_fd_sc_hd__buf_12
Xoutput88 net88 VGND VGND VPWR VPWR debug_reg3[30] sky130_fd_sc_hd__buf_8
Xoutput77 net77 VGND VGND VPWR VPWR debug_reg3[20] sky130_fd_sc_hd__buf_8
XFILLER_0_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput99 net99 VGND VGND VPWR VPWR instruction_debug[21] sky130_fd_sc_hd__buf_8
XFILLER_0_37_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1620_ net212 _0515_ _0516_ net4 VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1551_ net252 _0504_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1482_ net484 _0487_ _0489_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1818_ clknet_leaf_8_clk net279 VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_100_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold310 net134 VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1749_ clknet_leaf_9_clk _0066_ VGND VGND VPWR VPWR ex_mem_valid sky130_fd_sc_hd__dfxtp_1
Xhold321 net113 VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 _0562_ VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold343 register_file.write_data\[10\] VGND VGND VPWR VPWR net538 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0982_ dmem.address\[5\] _0619_ _0620_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_132_Right_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1603_ _0511_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1534_ net58 _0503_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1465_ _0452_ _0478_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1396_ _0440_ net330 net434 VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__nor3b_1
XTAP_TAPCELL_ROW_2_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold162 net53 VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 _0269_ VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold140 dmem.address\[20\] VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold184 _0204_ VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 _0177_ VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 net62 VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1250_ net326 _0308_ _0692_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__mux2_1
X_1181_ _0780_ _0792_ _0806_ _0607_ VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__a31o_1
XFILLER_0_87_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0965_ _0589_ _0591_ _0604_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0896_ register_file.write_data\[0\] _0538_ net141 _0535_ net543 VGND VGND VPWR VPWR
+ _0540_ sky130_fd_sc_hd__a32o_1
XFILLER_0_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1517_ net228 _0500_ _0501_ net288 VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__a22o_1
X_1448_ net451 _0467_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1379_ register_file.write_data\[31\] id_ex_rs2_data\[31\] _0833_ VGND VGND VPWR
+ VPWR _0429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1302_ _0345_ _0344_ _0357_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__a21oi_1
X_1233_ _0794_ _0291_ _0292_ _0837_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_88_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1164_ _0782_ _0790_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_74 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1095_ _0725_ _0726_ VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0948_ _0586_ _0588_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0879_ _0525_ net437 VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1920_ clknet_leaf_7_clk _0236_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_126_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1851_ clknet_leaf_8_clk net350 VGND VGND VPWR VPWR id_ex_rs2_data\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1782_ clknet_leaf_13_clk _0098_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1216_ _0773_ _0832_ _0838_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1147_ dmem.address\[16\] _0611_ VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1078_ _0707_ _0708_ _0710_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold22 _0223_ VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 register_file.write_data\[16\] VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 net80 VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 _0124_ VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 register_file.write_data\[20\] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 _0133_ VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold77 net36 VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 _0246_ VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 register_file.write_data\[1\] VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1001_ net139 _0638_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1903_ clknet_leaf_1_clk net209 VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_45_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1834_ clknet_leaf_0_clk net384 VGND VGND VPWR VPWR id_ex_rs2_data\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1765_ clknet_leaf_15_clk net332 VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_25_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1696_ clknet_leaf_3_clk _0013_ VGND VGND VPWR VPWR register_file.write_data\[12\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_0_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput34 net34 VGND VGND VPWR VPWR debug_reg2[10] sky130_fd_sc_hd__buf_8
Xoutput12 net12 VGND VGND VPWR VPWR debug_reg1[1] sky130_fd_sc_hd__buf_8
Xoutput23 net23 VGND VGND VPWR VPWR debug_reg1[2] sky130_fd_sc_hd__buf_8
Xoutput67 net67 VGND VGND VPWR VPWR debug_reg3[11] sky130_fd_sc_hd__buf_8
Xoutput56 net56 VGND VGND VPWR VPWR debug_reg2[30] sky130_fd_sc_hd__buf_8
Xoutput45 net45 VGND VGND VPWR VPWR debug_reg2[20] sky130_fd_sc_hd__buf_8
Xoutput89 net89 VGND VGND VPWR VPWR debug_reg3[31] sky130_fd_sc_hd__buf_8
Xoutput78 net78 VGND VGND VPWR VPWR debug_reg3[21] sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_8_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_113_Right_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1550_ net266 _0504_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1481_ _0452_ _0488_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_91_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1817_ clknet_leaf_8_clk net283 VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_100_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold300 id_ex_rs1_data\[26\] VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_68_Left_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold311 id_ex_immediate\[0\] VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1748_ clknet_leaf_9_clk _0065_ VGND VGND VPWR VPWR mem_wb_valid sky130_fd_sc_hd__dfxtp_2
XFILLER_0_102_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold322 _0472_ VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 net50 VGND VGND VPWR VPWR net539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 _0563_ VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1679_ net404 _0239_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_51_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_77_Left_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_86_Left_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0981_ _0532_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__buf_4
XFILLER_0_39_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1602_ net308 _0493_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__nor2_4
XFILLER_0_2_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1533_ net419 _0503_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__and2_1
X_1464_ net449 _0477_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1395_ reset net129 net499 net472 VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__or4_4
XFILLER_0_38_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold130 _0027_ VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 net52 VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 _0021_ VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold163 _0201_ VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 dmem.address\[18\] VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 _0148_ VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold196 net95 VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_21_clk net175 VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1180_ _0780_ _0792_ _0806_ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_12_clk net190 VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_8
X_0964_ _0586_ _0588_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0895_ net313 forwarding_unit.rs2_ex\[3\] forwarding_unit.rs2_ex\[0\] forwarding_unit.rs2_ex\[1\]
+ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1516_ net202 _0500_ _0501_ net232 VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1447_ _0522_ net467 _0467_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__nor3_1
X_1378_ _0413_ _0416_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_14_Left_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Left_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1301_ _0355_ _0356_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__or2b_1
X_1232_ dmem.address\[21\] _0835_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_1_clk net179 VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_88_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1163_ _0782_ _0790_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_32_Left_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1094_ _0719_ _0721_ _0724_ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__nand3_1
XFILLER_0_87_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0947_ net436 _0587_ _0532_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0878_ _0525_ net435 VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Left_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Left_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload0 clknet_1_1__leaf_clk VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__inv_8
XFILLER_0_123_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1850_ clknet_leaf_5_clk _0166_ VGND VGND VPWR VPWR id_ex_rs2_data\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1781_ clknet_leaf_13_clk net448 VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_127_Right_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1215_ _0773_ _0832_ _0838_ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__or3_1
XFILLER_0_79_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1146_ register_file.write_data\[16\] id_ex_rs2_data\[16\] _0609_ VGND VGND VPWR
+ VPWR _0774_ sky130_fd_sc_hd__mux2_1
X_1077_ net414 _0709_ _0532_ VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold23 register_file.write_data\[11\] VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 _0221_ VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 _0132_ VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 net68 VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 _0225_ VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold78 _0185_ VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 net38 VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 net31 VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1000_ _0603_ _0605_ _0622_ _0601_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_106_Left_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1902_ clknet_leaf_1_clk net221 VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_120_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1833_ clknet_leaf_21_clk _0149_ VGND VGND VPWR VPWR id_ex_rs2_data\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1764_ clknet_leaf_16_clk _0080_ VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1695_ clknet_leaf_3_clk _0012_ VGND VGND VPWR VPWR register_file.write_data\[11\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_40_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1129_ _0734_ _0746_ _0758_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_105_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput13 net13 VGND VGND VPWR VPWR debug_reg1[20] sky130_fd_sc_hd__buf_12
Xoutput24 net24 VGND VGND VPWR VPWR debug_reg1[30] sky130_fd_sc_hd__buf_8
Xoutput57 net57 VGND VGND VPWR VPWR debug_reg2[31] sky130_fd_sc_hd__buf_8
Xoutput46 net46 VGND VGND VPWR VPWR debug_reg2[21] sky130_fd_sc_hd__buf_8
Xoutput35 net35 VGND VGND VPWR VPWR debug_reg2[11] sky130_fd_sc_hd__buf_8
Xoutput79 net79 VGND VGND VPWR VPWR debug_reg3[22] sky130_fd_sc_hd__buf_8
Xoutput68 net68 VGND VGND VPWR VPWR debug_reg3[12] sky130_fd_sc_hd__buf_8
XFILLER_0_98_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1480_ net484 _0487_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1816_ clknet_leaf_9_clk net251 VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_100_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold301 _0061_ VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1747_ clknet_leaf_10_clk _0064_ VGND VGND VPWR VPWR dmem.address\[31\] sky130_fd_sc_hd__dfxtp_1
Xhold323 net110 VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 _0545_ VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 _0034_ VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold345 net122 VGND VGND VPWR VPWR net540 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1678_ net408 _0239_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0980_ register_file.write_data\[5\] id_ex_rs1_data\[5\] _0618_ VGND VGND VPWR VPWR
+ _0619_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1601_ net378 net314 _0507_ net57 VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1532_ net44 _0503_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__and2_1
X_1463_ _0564_ net427 _0477_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__nor3_1
XFILLER_0_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1394_ net131 net130 net471 net132 VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__or4_1
XFILLER_0_38_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold153 _0168_ VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 _0198_ VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 dmem.address\[22\] VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 net359 VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__clkbuf_4
Xhold175 dmem.address\[19\] VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 _0019_ VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 net97 VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold197 net88 VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0963_ net398 _0602_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0894_ net313 net308 net386 VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__o21a_2
XFILLER_0_55_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1515_ net216 _0500_ _0501_ net244 VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1446_ net518 net466 _0463_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__and3_1
X_1377_ _0411_ _0426_ _0427_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_108_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1300_ _0352_ _0354_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1231_ register_file.write_data\[21\] id_ex_rs2_data\[21\] _0833_ VGND VGND VPWR
+ VPWR _0291_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1162_ _0784_ _0789_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1093_ _0719_ _0721_ _0724_ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1995_ if_id_valid VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_31_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0946_ register_file.write_data\[3\] id_ex_rs1_data\[3\] _0528_ VGND VGND VPWR VPWR
+ _0587_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0877_ _0525_ net200 VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1429_ net134 _0453_ net502 VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_126_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload1 clknet_leaf_5_clk VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_19_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1780_ clknet_leaf_13_clk net465 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1214_ _0794_ _0834_ _0836_ _0837_ VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1145_ _0772_ VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__buf_2
XFILLER_0_94_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1076_ register_file.write_data\[11\] id_ex_rs1_data\[11\] _0528_ VGND VGND VPWR
+ VPWR _0709_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0929_ dmem.address\[2\] _0537_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold13 register_file.write_data\[14\] VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 _0121_ VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 dmem.address\[4\] VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 _0216_ VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 net43 VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 net37 VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 _0187_ VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_45 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1901_ clknet_leaf_1_clk net213 VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_45_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1832_ clknet_leaf_1_clk net369 VGND VGND VPWR VPWR id_ex_rs2_data\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_41_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1763_ clknet_leaf_15_clk _0079_ VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_40_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1694_ clknet_leaf_17_clk _0011_ VGND VGND VPWR VPWR register_file.write_data\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_40_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1128_ _0725_ _0744_ _0745_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1059_ net420 _0691_ _0692_ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput14 net14 VGND VGND VPWR VPWR debug_reg1[21] sky130_fd_sc_hd__buf_12
Xoutput25 net25 VGND VGND VPWR VPWR debug_reg1[31] sky130_fd_sc_hd__buf_8
XFILLER_0_113_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput47 net47 VGND VGND VPWR VPWR debug_reg2[22] sky130_fd_sc_hd__buf_8
Xoutput36 net36 VGND VGND VPWR VPWR debug_reg2[12] sky130_fd_sc_hd__buf_8
XFILLER_0_12_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput58 net58 VGND VGND VPWR VPWR debug_reg2[3] sky130_fd_sc_hd__buf_12
Xoutput69 net69 VGND VGND VPWR VPWR debug_reg3[13] sky130_fd_sc_hd__buf_8
XFILLER_0_11_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1815_ clknet_leaf_9_clk net249 VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_100_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold302 net127 VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1746_ clknet_leaf_10_clk _0063_ VGND VGND VPWR VPWR dmem.address\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold313 _0547_ VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 id_ex_rs1_data\[1\] VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold324 net11 VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold346 net119 VGND VGND VPWR VPWR net541 sky130_fd_sc_hd__dlygate4sd3_1
X_1677_ net490 _0239_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_125_Left_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1600_ net372 net314 _0507_ net56 VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1531_ net33 _0503_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__and2_1
X_1462_ net426 net117 _0473_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1393_ net105 net134 net106 VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_2_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold110 _0195_ VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold143 _0271_ VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 _0023_ VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 net46 VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1729_ clknet_leaf_17_clk _0046_ VGND VGND VPWR VPWR dmem.address\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold154 net51 VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 _0020_ VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 _0253_ VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold198 net89 VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 dmem.address\[14\] VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0962_ net397 _0600_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0893_ _0535_ net142 VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__nand2_2
XFILLER_0_15_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1514_ net214 _0500_ _0501_ net242 VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1445_ net110 _0463_ net466 VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__a21oi_1
X_1376_ _0412_ _0424_ _0425_ _0422_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_128_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1230_ _0284_ _0289_ _0290_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1161_ _0731_ _0783_ _0787_ _0788_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1092_ net438 _0556_ _0723_ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1994_ id_ex_valid VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__buf_1
XFILLER_0_27_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0945_ _0584_ net521 VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0876_ _0525_ net324 VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1428_ net505 _0453_ _0455_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__o21a_1
X_1359_ _0522_ _0409_ _0410_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_39_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_108_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload2 clknet_leaf_10_clk VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_80_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1213_ _0613_ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1144_ _0660_ _0706_ _0752_ _0765_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__or4_1
X_1075_ _0660_ _0687_ _0705_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0928_ id_ex_rs2_data\[2\] _0566_ _0568_ _0569_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__a211o_1
XFILLER_0_3_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0859_ _0000_ net414 VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold14 _0219_ VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 net73 VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 _0005_ VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 register_file.write_data\[13\] VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 _0192_ VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 net28 VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_66_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1900_ clknet_leaf_1_clk net219 VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__dfxtp_2
X_1831_ clknet_leaf_1_clk net367 VGND VGND VPWR VPWR id_ex_rs2_data\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_41_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1762_ clknet_leaf_19_clk _0078_ VGND VGND VPWR VPWR forwarding_unit.reg_write_wb
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1693_ clknet_leaf_19_clk _0010_ VGND VGND VPWR VPWR register_file.write_data\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Left_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1127_ _0754_ _0756_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_49_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1058_ _0620_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__buf_4
XFILLER_0_48_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Left_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput15 net15 VGND VGND VPWR VPWR debug_reg1[22] sky130_fd_sc_hd__buf_12
Xoutput48 net48 VGND VGND VPWR VPWR debug_reg2[23] sky130_fd_sc_hd__buf_8
Xoutput37 net37 VGND VGND VPWR VPWR debug_reg2[13] sky130_fd_sc_hd__buf_8
Xoutput26 net26 VGND VGND VPWR VPWR debug_reg1[3] sky130_fd_sc_hd__buf_8
XFILLER_0_12_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_47_Left_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput59 net59 VGND VGND VPWR VPWR debug_reg2[4] sky130_fd_sc_hd__buf_12
XFILLER_0_98_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_56_Left_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1814_ clknet_leaf_9_clk net287 VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_100_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1745_ clknet_leaf_10_clk _0062_ VGND VGND VPWR VPWR dmem.address\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_133_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold325 id_ex_immediate\[3\] VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 _0033_ VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold303 net106 VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__dlygate4sd3_1
X_1676_ net337 _0592_ net487 VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold336 _0560_ VGND VGND VPWR VPWR net531 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1530_ net140 VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__clkbuf_2
X_1461_ net426 _0473_ net117 VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1392_ net459 _0628_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_15_clk net192 VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_116_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold100 _0174_ VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 net20 VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 dmem.address\[23\] VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 net48 VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 _0194_ VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1728_ clknet_leaf_17_clk _0045_ VGND VGND VPWR VPWR dmem.address\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold177 register_file.write_data\[30\] VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 _0167_ VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold166 net2 VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__dlygate4sd3_1
X_1659_ _0517_ _0518_ net6 VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_113_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold199 net96 VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 net64 VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0961_ net397 _0600_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0892_ forwarding_unit.rd_mem\[0\] forwarding_unit.rs2_ex\[3\] forwarding_unit.rs2_ex\[0\]
+ forwarding_unit.rs2_ex\[1\] VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1513_ net206 _0500_ _0501_ net236 VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1444_ net514 _0463_ _0465_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_4_clk net188 VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_8
X_1375_ _0412_ _0422_ _0424_ _0425_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_128_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_122_Right_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1160_ _0757_ _0758_ _0769_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_88_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1091_ id_ex_rs1_data\[12\] _0558_ _0722_ _0620_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1993_ ex_mem_valid VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_31_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0944_ _0553_ _0572_ _0582_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0875_ _0525_ net421 VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Left_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1427_ net505 _0453_ _0564_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__a21oi_1
X_1358_ _0400_ _0398_ _0408_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_39_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1289_ _0339_ _0341_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__or2b_1
XFILLER_0_78_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload3 clknet_leaf_11_clk VGND VGND VPWR VPWR clkload3/Y sky130_fd_sc_hd__inv_12
XFILLER_0_18_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1212_ dmem.address\[20\] _0835_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_125_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1143_ _0770_ _0771_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__nor2_1
X_1074_ _0660_ _0706_ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0927_ register_file.write_data\[2\] _0538_ net141 VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0858_ _0000_ net420 VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold37 net75 VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 register_file.write_data\[10\] VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 _0218_ VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 _0126_ VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 net40 VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1830_ clknet_leaf_2_clk _0146_ VGND VGND VPWR VPWR id_ex_rs2_data\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1761_ clknet_leaf_19_clk _0077_ VGND VGND VPWR VPWR forwarding_unit.rd_mem\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1692_ clknet_leaf_19_clk _0009_ VGND VGND VPWR VPWR register_file.write_data\[8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_123_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1126_ net382 _0755_ _0620_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_105_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1057_ net538 id_ex_rs1_data\[10\] _0690_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1959_ clknet_leaf_18_clk _0275_ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput49 net49 VGND VGND VPWR VPWR debug_reg2[24] sky130_fd_sc_hd__buf_8
Xoutput38 net38 VGND VGND VPWR VPWR debug_reg2[14] sky130_fd_sc_hd__buf_8
XFILLER_0_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput27 net27 VGND VGND VPWR VPWR debug_reg1[4] sky130_fd_sc_hd__buf_8
Xoutput16 net16 VGND VGND VPWR VPWR debug_reg1[23] sky130_fd_sc_hd__buf_12
XFILLER_0_98_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_clk net169 VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1813_ clknet_leaf_9_clk net289 VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_100_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1744_ clknet_leaf_10_clk net496 VGND VGND VPWR VPWR dmem.address\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold315 id_reg_write VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 _0585_ VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold304 _0438_ VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1675_ net337 _0592_ net353 VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold337 _0035_ VGND VGND VPWR VPWR net532 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1109_ _0646_ _0720_ _0718_ _0737_ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_24_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Left_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1460_ net426 _0473_ _0475_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__o21a_1
X_1391_ net533 _0628_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold101 register_file.write_data\[8\] VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold123 net49 VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 _0024_ VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 _0196_ VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1727_ clknet_leaf_17_clk _0044_ VGND VGND VPWR VPWR dmem.address\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold156 register_file.write_data\[28\] VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 _0267_ VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 net3 VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__dlygate4sd3_1
X_1658_ _0517_ _0518_ net5 VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold178 _0203_ VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 _0150_ VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__dlygate4sd3_1
X_1589_ net202 _0509_ _0510_ net252 VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0960_ net230 _0599_ _0532_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0891_ forwarding_unit.rd_mem\[0\] forwarding_unit.rd_mem\[1\] net433 VGND VGND VPWR
+ VPWR _0535_ sky130_fd_sc_hd__o21a_1
XFILLER_0_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1512_ net204 _0500_ _0501_ net238 VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1443_ net514 _0463_ _0564_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1374_ _0405_ _0407_ _0400_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_74_Left_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_83_Left_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_92_Left_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1090_ register_file.write_data\[12\] _0618_ VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1992_ mem_wb_valid VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_7_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0943_ _0583_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__buf_2
XFILLER_0_15_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0874_ _0519_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__buf_1
Xclkload10 clknet_leaf_14_clk VGND VGND VPWR VPWR clkload10/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_55_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_578 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1426_ net471 net492 _0454_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__o21a_1
X_1357_ _0400_ _0398_ _0408_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__nor3b_1
XTAP_TAPCELL_ROW_39_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_52 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1288_ _0343_ _0344_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__nor2b_1
XFILLER_0_78_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload4 clknet_leaf_19_clk VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_18_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1211_ _0611_ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_125_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1142_ _0762_ _0761_ _0769_ _0607_ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1073_ _0687_ _0705_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0926_ _0530_ _0567_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0857_ _0000_ net425 VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold38 _0128_ VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold27 register_file.write_data\[23\] VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__dlygate4sd3_1
X_1409_ net330 net434 VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__xnor2_1
Xhold16 _0215_ VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 net74 VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1760_ clknet_leaf_18_clk net334 VGND VGND VPWR VPWR forwarding_unit.rd_mem\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_41_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1691_ clknet_leaf_0_clk net199 VGND VGND VPWR VPWR register_file.write_data\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_123_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1125_ register_file.write_data\[14\] id_ex_rs1_data\[14\] _0618_ VGND VGND VPWR
+ VPWR _0755_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1056_ _0618_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__buf_4
XFILLER_0_8_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1958_ clknet_leaf_19_clk _0274_ VGND VGND VPWR VPWR id_ex_immediate\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1889_ clknet_leaf_21_clk _0205_ VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__dfxtp_1
X_0909_ _0537_ _0549_ _0550_ _0551_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__a31o_1
XFILLER_0_16_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput39 net39 VGND VGND VPWR VPWR debug_reg2[15] sky130_fd_sc_hd__buf_8
Xoutput28 net28 VGND VGND VPWR VPWR debug_reg1[5] sky130_fd_sc_hd__buf_8
Xoutput17 net17 VGND VGND VPWR VPWR debug_reg1[24] sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_67_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_117_Right_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1812_ clknet_leaf_9_clk net233 VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1743_ clknet_leaf_11_clk _0060_ VGND VGND VPWR VPWR dmem.address\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold316 net122 VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__dlygate4sd3_1
X_1674_ net337 _0592_ net345 VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__and3_1
Xhold305 net131 VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold327 _0589_ VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 forwarding_unit.rd_mem\[0\] VGND VGND VPWR VPWR net533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1108_ _0660_ _0706_ _0738_ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__or3_1
XFILLER_0_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1039_ _0526_ _0541_ id_ex_rs2_data\[9\] VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_24_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_length12 net181 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_63_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_103_Left_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_112_Left_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1390_ _0525_ net413 VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_121_Left_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_130_Left_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_551 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold124 _0197_ VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 _0181_ VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold135 net128 VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 forwarding_unit.rd_wb\[1\] VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__dlygate4sd3_1
X_1726_ clknet_leaf_17_clk _0043_ VGND VGND VPWR VPWR dmem.address\[10\] sky130_fd_sc_hd__dfxtp_1
Xhold146 register_file.write_data\[29\] VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 _0137_ VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__dlygate4sd3_1
X_1657_ _0517_ _0518_ net365 VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__and3_1
Xhold168 net9 VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1588_ net216 _0509_ _0510_ net266 VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__a22o_1
Xhold179 dmem.address\[17\] VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0890_ net506 net395 VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1511_ net208 _0500_ _0501_ net234 VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1442_ net109 net416 _0464_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1373_ _0360_ _0362_ _0395_ _0396_ _0423_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__a311o_1
XFILLER_0_65_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1709_ clknet_leaf_5_clk _0026_ VGND VGND VPWR VPWR register_file.write_data\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1991_ net100 VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__buf_1
XFILLER_0_27_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0942_ _0553_ _0572_ _0582_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__or3_1
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0873_ _0524_ net430 VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload11 clknet_leaf_15_clk VGND VGND VPWR VPWR clkload11/Y sky130_fd_sc_hd__inv_8
XFILLER_0_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1425_ _0452_ _0453_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__nor2_1
X_1356_ _0405_ _0407_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_39_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1287_ _0329_ _0334_ _0342_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload5 clknet_leaf_20_clk VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__inv_6
XFILLER_0_61_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1210_ register_file.write_data\[20\] id_ex_rs2_data\[20\] _0833_ VGND VGND VPWR
+ VPWR _0834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1141_ _0762_ _0761_ _0769_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_125_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1072_ _0594_ _0703_ _0704_ _0613_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0925_ forwarding_unit.rd_mem\[0\] forwarding_unit.rs2_ex\[3\] forwarding_unit.rs2_ex\[0\]
+ forwarding_unit.rs2_ex\[1\] VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__or4b_1
XFILLER_0_125_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0856_ _0000_ net423 VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1408_ _0522_ net434 VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__nor2_1
Xhold17 register_file.write_data\[12\] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 _0228_ VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 net70 VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__dlygate4sd3_1
X_1339_ net351 id_ex_rs1_data\[28\] _0690_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1690_ clknet_leaf_0_clk net197 VGND VGND VPWR VPWR register_file.write_data\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_52_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1124_ _0739_ _0751_ _0753_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_49_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1055_ _0660_ _0687_ _0688_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_105_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1957_ clknet_leaf_19_clk _0273_ VGND VGND VPWR VPWR id_ex_immediate\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1888_ clknet_leaf_8_clk net379 VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0908_ ex_mem_alu_result\[1\] _0535_ net142 net395 VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput29 net29 VGND VGND VPWR VPWR debug_reg1[6] sky130_fd_sc_hd__buf_8
Xoutput18 net18 VGND VGND VPWR VPWR debug_reg1[25] sky130_fd_sc_hd__buf_8
XFILLER_0_11_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1811_ clknet_leaf_9_clk net245 VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1742_ clknet_leaf_11_clk _0059_ VGND VGND VPWR VPWR dmem.address\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold317 net119 VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__dlygate4sd3_1
X_1673_ net337 _0592_ net355 VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__and3_1
Xhold306 net23 VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold328 _0036_ VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 net103 VGND VGND VPWR VPWR net534 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_18_clk net185 VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1107_ _0718_ _0737_ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__nand2_1
X_1038_ register_file.write_data\[9\] _0538_ net542 VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_length24 net193 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__buf_1
XFILLER_0_118_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1725_ clknet_leaf_17_clk _0042_ VGND VGND VPWR VPWR dmem.address\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold125 net45 VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 _0511_ VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__clkbuf_4
Xhold103 net32 VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 _0138_ VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 net24 VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk net181 VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold136 _0444_ VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__dlygate4sd3_1
X_1656_ _0517_ _0518_ net362 VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_113_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1587_ net214 _0509_ _0510_ net268 VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold169 net13 VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1510_ net220 _0500_ _0501_ net246 VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1441_ _0452_ _0463_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1372_ _0394_ _0408_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_128_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1708_ clknet_leaf_5_clk _0025_ VGND VGND VPWR VPWR register_file.write_data\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1639_ net378 net309 _0513_ net487 VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_70_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1990_ net99 VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__buf_1
XFILLER_0_27_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0941_ _0543_ net520 _0580_ _0581_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_31_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0872_ _0524_ net328 VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload12 clknet_leaf_16_clk VGND VGND VPWR VPWR clkload12/Y sky130_fd_sc_hd__inv_8
XFILLER_0_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1424_ net500 net471 net491 _0446_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__and4_1
X_1355_ net437 _0406_ _0692_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1286_ _0329_ _0334_ _0342_ _0521_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_39_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload6 clknet_leaf_21_clk VGND VGND VPWR VPWR clkload6/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_116_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1140_ _0766_ _0768_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_125_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1071_ dmem.address\[11\] _0611_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0924_ _0538_ net141 VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__nand2_2
XFILLER_0_28_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0855_ _0000_ net198 VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold29 register_file.write_data\[22\] VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__dlygate4sd3_1
X_1407_ net433 _0628_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__and2_1
Xhold18 _0217_ VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__dlygate4sd3_1
X_1338_ _0378_ _0390_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1269_ _0325_ _0326_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_89_Left_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_98_Left_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_49 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1123_ _0660_ _0706_ _0752_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_49_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1054_ _0660_ _0683_ _0686_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_105_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1956_ clknet_leaf_19_clk _0272_ VGND VGND VPWR VPWR id_ex_immediate\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0907_ _0538_ net141 id_ex_rs2_data\[1\] VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__a21o_1
X_1887_ clknet_leaf_8_clk net373 VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_131_Right_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput19 net19 VGND VGND VPWR VPWR debug_reg1[26] sky130_fd_sc_hd__buf_8
XFILLER_0_101_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1810_ clknet_leaf_9_clk net243 VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1741_ clknet_leaf_5_clk _0058_ VGND VGND VPWR VPWR dmem.address\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1672_ net337 _0592_ net339 VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold307 net105 VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold318 _0101_ VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 net15 VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1106_ _0594_ _0735_ _0736_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1037_ _0584_ _0615_ _0645_ _0664_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__or4_1
XFILLER_0_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_length14 net183 VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_75_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1939_ clknet_leaf_3_clk _0255_ VGND VGND VPWR VPWR id_ex_rs1_data\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Left_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1724_ clknet_leaf_17_clk _0041_ VGND VGND VPWR VPWR dmem.address\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold115 _0229_ VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 _0193_ VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 _0249_ VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold148 net54 VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 _0270_ VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold137 _0081_ VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__dlygate4sd3_1
X_1655_ _0519_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_44_Left_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1586_ net206 _0509_ _0510_ net254 VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_53_Left_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Left_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1440_ net109 net416 VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__and2_1
X_1371_ _0420_ _0421_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_128_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1707_ clknet_leaf_5_clk net329 VGND VGND VPWR VPWR register_file.write_data\[23\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_14_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1638_ net372 net309 _0513_ net353 VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1569_ net294 _0506_ _0508_ net44 VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_70_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Left_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_109_Left_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0940_ dmem.address\[3\] _0535_ net142 net395 VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0871_ _0524_ net326 VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_11_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload13 clknet_leaf_17_clk VGND VGND VPWR VPWR clkload13/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_51_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1423_ _0521_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_118_Left_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1354_ net536 id_ex_rs1_data\[29\] _0690_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__mux2_1
X_1285_ _0339_ _0341_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_39_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_127_Left_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload7 clknet_leaf_4_clk VGND VGND VPWR VPWR clkload7/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1070_ register_file.write_data\[11\] id_ex_rs2_data\[11\] _0609_ VGND VGND VPWR
+ VPWR _0703_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_112_Right_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0923_ _0546_ net528 _0565_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__o21a_1
XFILLER_0_28_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0854_ _0000_ net196 VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1406_ net441 _0628_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__and2_1
Xhold19 register_file.write_data\[17\] VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__dlygate4sd3_1
X_1337_ _0794_ _0388_ _0389_ _0837_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1268_ _0310_ _0316_ _0324_ _0607_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1199_ dmem.address\[19\] _0611_ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1122_ _0738_ _0751_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_79 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1053_ _0683_ _0686_ VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_49_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1955_ clknet_leaf_8_clk net338 VGND VGND VPWR VPWR id_ex_rs1_data\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_64_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0906_ register_file.write_data\[1\] _0526_ _0541_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__or3_1
XFILLER_0_22_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1886_ clknet_leaf_8_clk net344 VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1740_ clknet_leaf_5_clk _0057_ VGND VGND VPWR VPWR dmem.address\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1671_ net337 _0592_ net409 VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold308 _0456_ VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold319 net110 VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1105_ dmem.address\[13\] _0611_ _0613_ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__o21a_1
XFILLER_0_76_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1036_ _0665_ _0667_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_length26 net195 VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__buf_1
X_1938_ clknet_leaf_3_clk _0254_ VGND VGND VPWR VPWR id_ex_rs1_data\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_118_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1869_ clknet_leaf_2_clk net273 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1723_ clknet_leaf_19_clk _0040_ VGND VGND VPWR VPWR dmem.address\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold116 net18 VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold105 register_file.write_data\[0\] VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 _0202_ VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 dmem.address\[21\] VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 id_ex_rd_addr\[0\] VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__dlygate4sd3_1
X_1654_ net337 VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_110_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1585_ net204 _0509_ _0510_ net256 VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1019_ _0654_ _0655_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1370_ _0419_ _0417_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_128_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1706_ clknet_leaf_5_clk net327 VGND VGND VPWR VPWR register_file.write_data\[22\]
+ sky130_fd_sc_hd__dfxtp_2
X_1637_ net341 net309 _0513_ net345 VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1568_ net300 _0506_ _0508_ net33 VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__a22o_1
X_1499_ register_file.write_data\[4\] _0497_ _0499_ net454 VGND VGND VPWR VPWR _0113_
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_126_Right_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0870_ _0524_ net322 VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_11_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload14 clknet_leaf_18_clk VGND VGND VPWR VPWR clkload14/Y sky130_fd_sc_hd__inv_8
XFILLER_0_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1422_ _0522_ _0450_ net492 VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__nor3_1
XFILLER_0_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1353_ _0401_ _0404_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__xnor2_1
X_1284_ net430 _0340_ _0692_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload8 clknet_leaf_12_clk VGND VGND VPWR VPWR clkload8/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_61_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0999_ _0635_ _0636_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_125_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0922_ _0546_ _0563_ _0564_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0853_ _0000_ net432 VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1405_ _0442_ net333 VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__and2_1
X_1336_ dmem.address\[28\] _0835_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1267_ _0310_ _0316_ _0324_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_69_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1198_ register_file.write_data\[19\] id_ex_rs2_data\[19\] _0609_ VGND VGND VPWR
+ VPWR _0823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1121_ _0594_ _0749_ _0750_ _0613_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1052_ _0594_ _0684_ _0685_ _0613_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_49_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1954_ clknet_leaf_8_clk net354 VGND VGND VPWR VPWR id_ex_rs1_data\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_64_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0905_ _0543_ net526 VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1885_ clknet_leaf_8_clk net358 VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1319_ _0372_ _0373_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_530 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1670_ net337 _0592_ net311 VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_133_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold309 _0087_ VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1104_ register_file.write_data\[13\] id_ex_rs2_data\[13\] _0609_ VGND VGND VPWR
+ VPWR _0735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1035_ _0628_ _0669_ _0670_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_length16 clknet_1_0__leaf_clk VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__buf_1
XFILLER_0_33_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_length27 clknet_1_1__leaf_clk VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__buf_1
X_1937_ clknet_leaf_0_clk net360 VGND VGND VPWR VPWR id_ex_rs1_data\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_118_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1868_ clknet_leaf_2_clk net277 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1799_ clknet_leaf_7_clk _0115_ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_77_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1722_ clknet_leaf_19_clk _0039_ VGND VGND VPWR VPWR dmem.address\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold117 _0230_ VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1653_ _0441_ _0411_ net361 VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__and3_1
Xhold106 _0173_ VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold128 _0022_ VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 _0076_ VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1584_ net208 _0509_ _0510_ net262 VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_113_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_107_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1018_ _0635_ _0641_ _0653_ _0607_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1705_ clknet_leaf_5_clk net323 VGND VGND VPWR VPWR register_file.write_data\[21\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1636_ net351 net309 _0513_ net355 VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_74_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1567_ _0507_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1498_ net292 _0497_ _0499_ net443 VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1421_ net131 net491 _0446_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_110_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1352_ _0794_ _0402_ _0403_ _0837_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__o211a_1
X_1283_ register_file.write_data\[24\] id_ex_rs1_data\[24\] _0690_ VGND VGND VPWR
+ VPWR _0340_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload9 clknet_leaf_13_clk VGND VGND VPWR VPWR clkload9/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_61_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0998_ _0634_ _0632_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__or2b_1
XFILLER_0_14_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1619_ _0513_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_59_Left_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0921_ _0521_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_44_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0852_ _0000_ net230 VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1404_ _0442_ net431 VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__and2_1
X_1335_ register_file.write_data\[28\] id_ex_rs2_data\[28\] _0833_ VGND VGND VPWR
+ VPWR _0388_ sky130_fd_sc_hd__mux2_1
X_1266_ _0321_ _0323_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_69_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1197_ _0819_ _0821_ _0822_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_82_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_67_Left_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Left_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1120_ dmem.address\[14\] _0611_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1051_ dmem.address\[10\] _0611_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_49_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1953_ clknet_leaf_8_clk net346 VGND VGND VPWR VPWR id_ex_rs1_data\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1884_ clknet_leaf_7_clk _0200_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dfxtp_1
X_0904_ _0546_ net508 _0522_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1318_ _0371_ _0360_ _0362_ _0607_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__a31o_1
X_1249_ register_file.write_data\[22\] id_ex_rs1_data\[22\] _0690_ VGND VGND VPWR
+ VPWR _0308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1103_ _0628_ _0733_ _0734_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_66_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1034_ _0658_ _0668_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1936_ clknet_leaf_0_clk _0252_ VGND VGND VPWR VPWR id_ex_rs1_data\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1867_ clknet_leaf_2_clk net271 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1798_ clknet_leaf_7_clk _0114_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_77_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1721_ clknet_leaf_0_clk net400 VGND VGND VPWR VPWR dmem.address\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1652_ _0441_ _0411_ net298 VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__and3_1
Xhold107 register_file.write_data\[9\] VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold129 dmem.address\[26\] VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold118 forwarding_unit.rd_wb\[0\] VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1583_ net220 _0509_ _0510_ net274 VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_13_Left_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1017_ _0635_ _0641_ _0653_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_22_Left_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1919_ clknet_leaf_7_clk _0235_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_60_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_31_Left_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Left_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1704_ clknet_leaf_5_clk net336 VGND VGND VPWR VPWR register_file.write_data\[20\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1635_ net494 net309 _0513_ net339 VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_74_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1566_ _0521_ net314 VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__nor2_4
XFILLER_0_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1497_ net290 _0497_ _0499_ net445 VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1420_ net500 _0446_ net491 VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1351_ dmem.address\[29\] _0835_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_56_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1282_ _0335_ _0338_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0997_ _0632_ _0634_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__or2b_1
XFILLER_0_131_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1618_ _0511_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1549_ net268 _0504_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_87_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold290 _0106_ VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_125_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0920_ _0561_ net527 VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_44_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0851_ _0000_ net436 VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1403_ _0519_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1334_ _0385_ _0386_ _0387_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__o21a_1
X_1265_ net328 _0322_ _0692_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1196_ _0819_ _0821_ _0592_ VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_82_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1050_ register_file.write_data\[10\] id_ex_rs2_data\[10\] _0609_ VGND VGND VPWR
+ VPWR _0684_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1952_ clknet_leaf_8_clk net356 VGND VGND VPWR VPWR id_ex_rs1_data\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_64_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1883_ clknet_leaf_7_clk _0199_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0903_ net507 _0533_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__or2b_1
XFILLER_0_43_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1317_ _0360_ _0362_ _0371_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1248_ _0295_ _0306_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__xor2_2
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1179_ _0804_ _0805_ VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__or2b_1
XFILLER_0_93_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1102_ _0727_ _0732_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1033_ _0658_ _0668_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1935_ clknet_leaf_0_clk _0251_ VGND VGND VPWR VPWR id_ex_rs1_data\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_length18 net188 VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__buf_1
XFILLER_0_133_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1866_ clknet_leaf_2_clk net303 VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1797_ clknet_leaf_7_clk _0113_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_95_Left_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_121_Right_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1720_ clknet_leaf_20_clk _0037_ VGND VGND VPWR VPWR dmem.address\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold108 _0182_ VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__dlygate4sd3_1
X_1651_ _0441_ _0411_ net284 VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__and3_1
Xhold119 _0505_ VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__clkbuf_4
X_1582_ net212 _0509_ _0510_ net272 VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_72_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1016_ _0651_ _0652_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1918_ clknet_leaf_7_clk _0234_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_8_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1849_ clknet_leaf_5_clk _0165_ VGND VGND VPWR VPWR id_ex_rs2_data\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_20_clk net175 VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_clk net183 VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1703_ clknet_leaf_3_clk net371 VGND VGND VPWR VPWR register_file.write_data\[19\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_30_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1634_ net280 net309 _0513_ net409 VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_74_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1565_ net314 VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__clkbuf_4
X_1496_ net294 _0497_ _0499_ net444 VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1350_ register_file.write_data\[29\] id_ex_rs2_data\[29\] _0833_ VGND VGND VPWR
+ VPWR _0402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1281_ _0794_ _0336_ _0337_ _0837_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_0_clk net179 VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_19_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0996_ net196 _0633_ _0620_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1617_ net218 _0512_ _0514_ net3 VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1548_ net254 _0504_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__and2_1
X_1479_ _0564_ net475 _0487_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_87_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold280 _0486_ VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 net26 VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_22 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0850_ _0000_ net422 VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1402_ _0525_ net534 VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__and2_1
X_1333_ _0385_ _0386_ _0564_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__a21oi_1
X_1264_ register_file.write_data\[23\] id_ex_rs1_data\[23\] _0690_ VGND VGND VPWR
+ VPWR _0322_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1195_ _0782_ _0790_ _0806_ _0820_ VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__o31a_1
XFILLER_0_36_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0979_ _0528_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_131_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_115_Left_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_124_Left_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_length6 clknet_0_clk VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_29_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1951_ clknet_leaf_8_clk net340 VGND VGND VPWR VPWR id_ex_rs1_data\[27\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_64_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1882_ clknet_leaf_6_clk net315 VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0902_ _0533_ _0545_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__or2b_1
XFILLER_0_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_133_Left_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1316_ _0369_ _0370_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__or2b_1
XFILLER_0_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1247_ _0794_ _0304_ _0305_ _0837_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__o211a_1
X_1178_ _0799_ _0800_ _0803_ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1101_ _0727_ _0732_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1032_ _0665_ _0667_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1934_ clknet_leaf_0_clk _0250_ VGND VGND VPWR VPWR id_ex_rs1_data\[10\] sky130_fd_sc_hd__dfxtp_1
Xmax_length19 net188 VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1865_ clknet_leaf_2_clk net297 VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1796_ clknet_leaf_7_clk _0112_ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1650_ _0441_ _0411_ net258 VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold109 net47 VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__dlygate4sd3_1
X_1581_ _0507_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1015_ _0646_ _0647_ _0650_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__or3_1
XFILLER_0_49_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1917_ clknet_leaf_7_clk _0233_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_71_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1848_ clknet_leaf_6_clk _0164_ VGND VGND VPWR VPWR id_ex_rs2_data\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1779_ clknet_leaf_13_clk _0095_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_9_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1702_ clknet_leaf_3_clk net381 VGND VGND VPWR VPWR register_file.write_data\[18\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_5_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1633_ net278 net309 _0513_ net311 VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_74_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1564_ net313 _0493_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__nor2_4
X_1495_ net300 _0497_ _0499_ net442 VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1280_ dmem.address\[24\] _0835_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0995_ register_file.write_data\[6\] id_ex_rs1_data\[6\] _0618_ VGND VGND VPWR VPWR
+ _0633_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1616_ net210 _0512_ _0514_ net2 VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1547_ net256 _0504_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__and2_1
X_1478_ net540 net474 _0483_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Left_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_28_Left_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold270 _0096_ VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold281 _0105_ VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 net25 VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_37_Left_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Left_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_116_Right_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1401_ _0525_ net404 VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__and2_1
X_1332_ _0369_ _0372_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__or2_1
X_1263_ _0317_ _0320_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1194_ _0780_ _0804_ _0805_ VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__o21a_1
XFILLER_0_36_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0978_ _0584_ net396 _0614_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__o21a_1
XFILLER_0_131_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1950_ clknet_leaf_5_clk _0266_ VGND VGND VPWR VPWR id_ex_rs1_data\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_64_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1881_ clknet_leaf_6_clk net319 VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0901_ _0534_ _0544_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1315_ _0366_ _0368_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1246_ dmem.address\[22\] _0835_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__or2_1
X_1177_ _0799_ _0800_ _0803_ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1100_ _0658_ _0728_ _0731_ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1031_ net423 _0666_ _0620_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1933_ clknet_leaf_0_clk net299 VGND VGND VPWR VPWR id_ex_rs1_data\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1864_ clknet_leaf_2_clk _0180_ VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1795_ clknet_leaf_7_clk _0111_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1229_ _0284_ _0289_ _0519_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1580_ net314 VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1014_ _0648_ _0650_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1916_ clknet_leaf_7_clk _0232_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_72_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1847_ clknet_leaf_6_clk _0163_ VGND VGND VPWR VPWR id_ex_rs2_data\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1778_ clknet_leaf_13_clk net452 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_9_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1701_ clknet_leaf_3_clk net375 VGND VGND VPWR VPWR register_file.write_data\[17\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_26_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1632_ net282 net309 _0513_ net17 VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1563_ net407 net140 VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_74_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1494_ _0498_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0994_ _0616_ _0631_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1615_ net302 _0512_ _0514_ net298 VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1546_ net262 _0504_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__and2_1
X_1477_ net122 _0483_ net474 VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_87_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold260 net121 VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 net111 VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 net27 VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 net60 VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_125_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1400_ _0525_ net408 VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__and2_1
X_1331_ _0383_ _0384_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__and2b_1
X_1262_ _0794_ _0318_ _0319_ _0837_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1193_ _0817_ _0818_ VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_82_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0977_ _0584_ _0615_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1529_ net100 net404 _0071_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0900_ net424 _0537_ _0540_ _0542_ _0543_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__o221a_1
XFILLER_0_113_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1880_ clknet_leaf_6_clk net307 VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1314_ _0366_ _0368_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__and2_1
X_1245_ register_file.write_data\[22\] id_ex_rs2_data\[22\] _0833_ VGND VGND VPWR
+ VPWR _0304_ sky130_fd_sc_hd__mux2_1
X_1176_ net374 _0556_ _0802_ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_48_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_65_Left_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1030_ register_file.write_data\[8\] id_ex_rs1_data\[8\] _0618_ VGND VGND VPWR VPWR
+ _0666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1932_ clknet_leaf_0_clk net285 VGND VGND VPWR VPWR id_ex_rs1_data\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1863_ clknet_leaf_2_clk _0179_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1794_ clknet_leaf_7_clk _0110_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1228_ _0790_ _0285_ _0288_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1159_ _0762_ _0785_ _0786_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_73_Left_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_82_Left_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_91_Left_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1013_ net198 _0649_ _0532_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1915_ clknet_leaf_7_clk _0231_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_60_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_14_clk net193 VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_127_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1846_ clknet_leaf_6_clk _0162_ VGND VGND VPWR VPWR id_ex_rs2_data\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1777_ clknet_leaf_13_clk net468 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1700_ clknet_leaf_3_clk net377 VGND VGND VPWR VPWR register_file.write_data\[16\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1631_ net222 _0515_ _0516_ net16 VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1562_ net406 net140 VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_74_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1493_ _0521_ _0496_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__nor2_4
XFILLER_0_10_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_3_clk net186 VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1829_ clknet_leaf_0_clk _0145_ VGND VGND VPWR VPWR id_ex_rs2_data\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0993_ _0594_ _0629_ _0630_ _0543_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1614_ net296 _0512_ _0514_ net284 VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__a22o_1
X_1545_ net274 _0504_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__and2_1
X_1476_ net511 _0483_ _0485_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__o21a_1
XFILLER_0_66_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold261 _0103_ VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__dlygate4sd3_1
Xhold250 net87 VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold272 _0466_ VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 net12 VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 _0178_ VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_130_Right_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1330_ _0378_ _0379_ _0382_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__nand3_1
X_1261_ dmem.address\[23\] _0835_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1192_ _0813_ _0814_ _0816_ VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__nor3_1
XFILLER_0_36_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0976_ net396 _0614_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__or2_2
XFILLER_0_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1528_ net378 _0496_ _0498_ net393 VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_93_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1459_ net426 _0473_ _0452_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_102_Left_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1313_ net324 _0367_ _0692_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__mux2_1
X_1244_ _0522_ _0303_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1175_ id_ex_rs1_data\[17\] _0558_ _0801_ _0620_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_48_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_111_Left_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0959_ register_file.write_data\[4\] id_ex_rs1_data\[4\] _0528_ VGND VGND VPWR VPWR
+ _0599_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_120_Left_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput130 net130 VGND VGND VPWR VPWR pc_current[5] sky130_fd_sc_hd__buf_8
XFILLER_0_30_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1931_ clknet_leaf_0_clk net259 VGND VGND VPWR VPWR id_ex_rs1_data\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1862_ clknet_leaf_2_clk net489 VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1793_ clknet_leaf_7_clk _0109_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1227_ _0819_ _0820_ _0829_ _0286_ _0287_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__o32ai_4
XFILLER_0_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1158_ _0766_ _0768_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1089_ _0646_ _0720_ _0718_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1012_ register_file.write_data\[7\] id_ex_rs1_data\[7\] _0528_ VGND VGND VPWR VPWR
+ _0649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1914_ clknet_leaf_6_clk net312 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_72_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1845_ clknet_leaf_6_clk _0161_ VGND VGND VPWR VPWR id_ex_rs2_data\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1776_ clknet_leaf_13_clk net515 VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1630_ net224 _0515_ _0516_ net15 VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1561_ net343 net140 VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_74_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1492_ _0496_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1828_ clknet_leaf_21_clk _0144_ VGND VGND VPWR VPWR id_ex_rs2_data\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_111_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1759_ clknet_leaf_9_clk _0000_ VGND VGND VPWR VPWR if_id_valid sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0992_ dmem.address\[6\] _0537_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1613_ register_file.write_data\[7\] _0512_ _0514_ net258 VGND VGND VPWR VPWR _0212_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1544_ net272 _0504_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1475_ net511 _0483_ _0452_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold240 dmem.address\[28\] VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 net94 VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 net107 VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 net126 VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 _0093_ VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 net99 VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1260_ register_file.write_data\[23\] id_ex_rs2_data\[23\] _0833_ VGND VGND VPWR
+ VPWR _0318_ sky130_fd_sc_hd__mux2_1
X_1191_ _0813_ _0814_ _0816_ VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__o21a_1
XFILLER_0_127_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_69_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0975_ _0594_ _0610_ _0612_ _0613_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1527_ net372 _0496_ _0498_ net392 VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_93_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1458_ net447 _0472_ _0474_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1389_ _0525_ net412 VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_124_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1312_ net410 net495 _0690_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1243_ _0301_ _0302_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1174_ register_file.write_data\[17\] _0618_ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_48_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0958_ _0584_ net396 VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_95_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0889_ net424 _0529_ _0532_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput120 net120 VGND VGND VPWR VPWR pc_current[25] sky130_fd_sc_hd__buf_8
Xoutput131 net131 VGND VGND VPWR VPWR pc_current[6] sky130_fd_sc_hd__buf_8
XFILLER_0_11_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1930_ clknet_leaf_0_clk net261 VGND VGND VPWR VPWR id_ex_rs1_data\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1861_ clknet_leaf_1_clk net390 VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_127_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1792_ clknet_leaf_12_clk _0108_ VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_clk net173 VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_1226_ _0826_ _0828_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1157_ _0766_ _0768_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1088_ _0687_ _0705_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_132_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_125_Right_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1011_ _0646_ _0647_ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1913_ clknet_leaf_6_clk net310 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_72_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1844_ clknet_leaf_6_clk _0160_ VGND VGND VPWR VPWR id_ex_rs2_data\[19\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_7_Left_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1775_ clknet_leaf_13_clk net417 VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1209_ _0609_ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__buf_4
XFILLER_0_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1560_ net357 net140 VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_74_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1491_ _0495_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1827_ clknet_leaf_0_clk _0143_ VGND VGND VPWR VPWR id_ex_rs2_data\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1758_ clknet_leaf_9_clk _0075_ VGND VGND VPWR VPWR id_ex_valid sky130_fd_sc_hd__dfxtp_1
Xmax_cap141 _0539_ VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_2
X_1689_ clknet_leaf_0_clk _0006_ VGND VGND VPWR VPWR register_file.write_data\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_127_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_79_Left_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_88_Left_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0991_ register_file.write_data\[6\] id_ex_rs2_data\[6\] _0566_ VGND VGND VPWR VPWR
+ _0629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1612_ register_file.write_data\[6\] _0512_ _0514_ net260 VGND VGND VPWR VPWR _0211_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_97_Left_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1543_ net140 VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1474_ net455 _0482_ _0484_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold252 net115 VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 dmem.address\[3\] VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold230 dmem.address\[9\] VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold285 _0107_ VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 net84 VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 net132 VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 _0461_ VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1190_ net380 _0815_ _0620_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0974_ _0543_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1526_ net341 _0496_ _0498_ net86 VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1457_ _0452_ _0473_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__nor2_1
X_1388_ _0436_ _0437_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_124_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_48 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1311_ _0350_ _0365_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__xnor2_1
X_1242_ _0284_ _0289_ _0281_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1173_ _0773_ _0776_ _0797_ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_87_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_25_Left_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0957_ _0594_ _0595_ _0596_ _0543_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput110 net110 VGND VGND VPWR VPWR pc_current[15] sky130_fd_sc_hd__buf_8
X_0888_ _0531_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput121 net121 VGND VGND VPWR VPWR pc_current[26] sky130_fd_sc_hd__buf_8
XFILLER_0_11_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput132 net132 VGND VGND VPWR VPWR pc_current[7] sky130_fd_sc_hd__buf_8
XFILLER_0_112_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1509_ net212 _0500_ _0501_ net240 VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_34_Left_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_106_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Left_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_52_Left_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Left_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1860_ clknet_leaf_1_clk net293 VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_126_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1791_ clknet_leaf_12_clk net480 VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1225_ _0826_ _0828_ _0817_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1156_ _0658_ _0728_ _0783_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__or3_1
XFILLER_0_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_17_clk net187 VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_8
X_1087_ _0660_ _0706_ _0718_ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__or3b_1
XFILLER_0_118_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1989_ net97 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__buf_1
XFILLER_0_16_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1010_ _0584_ _0615_ _0631_ _0644_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__o31a_1
XFILLER_0_44_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1912_ clknet_leaf_1_clk net223 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_121_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1843_ clknet_leaf_6_clk _0159_ VGND VGND VPWR VPWR id_ex_rs2_data\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1774_ clknet_leaf_14_clk _0090_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_6_clk net180 VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_108_Left_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1208_ _0812_ _0825_ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__or2_2
X_1139_ net385 _0767_ _0620_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_117_Left_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_126_Left_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1490_ net313 net308 _0494_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__and3_1
Xhold1 dmem.address\[6\] VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_85_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1826_ clknet_leaf_21_clk _0142_ VGND VGND VPWR VPWR id_ex_rs2_data\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1757_ clknet_leaf_19_clk _0074_ VGND VGND VPWR VPWR id_ex_rd_addr\[0\] sky130_fd_sc_hd__dfxtp_1
Xmax_cap142 net543 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__buf_1
XFILLER_0_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1688_ clknet_leaf_0_clk net231 VGND VGND VPWR VPWR register_file.write_data\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_111_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0990_ _0519_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__buf_1
XFILLER_0_26_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1611_ register_file.write_data\[5\] _0512_ _0514_ net264 VGND VGND VPWR VPWR _0210_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1542_ net276 _0503_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__and2_1
X_1473_ _0452_ _0483_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_558 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1809_ clknet_leaf_8_clk net237 VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold220 net108 VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold242 dmem.address\[29\] VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 net116 VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 _0097_ VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold275 _0136_ VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 forwarding_unit.rd_mem\[1\] VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 register_file.write_data\[7\] VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 _0451_ VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0973_ dmem.address\[5\] _0611_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1525_ net351 _0496_ _0498_ net85 VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_93_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1456_ net447 net517 VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__and2_1
X_1387_ _0420_ _0427_ _0435_ _0607_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1310_ _0794_ _0363_ _0364_ _0837_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__o211a_1
X_1241_ _0299_ _0300_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_47_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1172_ _0793_ _0798_ VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0956_ net230 _0537_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_95_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput100 net100 VGND VGND VPWR VPWR instruction_debug[22] sky130_fd_sc_hd__buf_8
X_0887_ _0530_ net459 forwarding_unit.rs1_ex\[0\] VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__or3b_1
Xoutput122 net122 VGND VGND VPWR VPWR pc_current[27] sky130_fd_sc_hd__buf_8
XFILLER_0_112_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput111 net111 VGND VGND VPWR VPWR pc_current[16] sky130_fd_sc_hd__buf_8
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput133 net133 VGND VGND VPWR VPWR pc_current[8] sky130_fd_sc_hd__buf_8
XFILLER_0_11_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1508_ _0498_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1439_ _0522_ net458 net416 VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__nor3_1
XFILLER_0_97_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1790_ clknet_leaf_12_clk net485 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1224_ _0782_ _0806_ _0819_ _0829_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__or4_1
XFILLER_0_79_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1155_ _0727_ _0746_ _0757_ _0769_ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__or4_1
X_1086_ _0594_ _0716_ _0717_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_87_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_74 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0939_ register_file.write_data\[3\] _0566_ _0537_ _0579_ VGND VGND VPWR VPWR _0580_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1911_ clknet_leaf_1_clk net225 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1842_ clknet_leaf_2_clk _0158_ VGND VGND VPWR VPWR id_ex_rs2_data\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1773_ clknet_leaf_14_clk _0089_ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1207_ _0829_ _0830_ _0831_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__o21a_1
XFILLER_0_95_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1138_ register_file.write_data\[15\] id_ex_rs1_data\[15\] _0618_ VGND VGND VPWR
+ VPWR _0767_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1069_ _0628_ _0701_ _0702_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_36_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2 _0007_ VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1825_ clknet_leaf_21_clk _0141_ VGND VGND VPWR VPWR id_ex_rs2_data\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1756_ clknet_leaf_19_clk _0073_ VGND VGND VPWR VPWR forwarding_unit.rs2_ex\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1687_ clknet_leaf_20_clk _0004_ VGND VGND VPWR VPWR register_file.write_data\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_0_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1610_ register_file.write_data\[4\] _0512_ _0514_ net477 VGND VGND VPWR VPWR _0209_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1541_ net270 _0503_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__and2_1
X_1472_ net455 _0482_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1808_ clknet_leaf_9_clk net239 VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold210 _0502_ VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 _0476_ VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__dlygate4sd3_1
X_1739_ clknet_leaf_4_clk _0056_ VGND VGND VPWR VPWR dmem.address\[23\] sky130_fd_sc_hd__dfxtp_1
Xhold221 _0462_ VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold243 dmem.address\[12\] VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold265 net120 VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 net118 VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 register_file.write_data\[6\] VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 net133 VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold298 _0085_ VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0972_ _0537_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_43_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1524_ register_file.write_data\[27\] _0496_ _0498_ net469 VGND VGND VPWR VPWR _0136_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1455_ _0522_ net464 _0472_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__nor3_1
X_1386_ _0420_ _0427_ _0435_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1240_ _0295_ _0296_ _0298_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__or3_1
X_1171_ _0776_ _0797_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_120_Right_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0955_ register_file.write_data\[4\] id_ex_rs2_data\[4\] _0566_ VGND VGND VPWR VPWR
+ _0595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0886_ forwarding_unit.rd_mem\[0\] forwarding_unit.rd_mem\[1\] forwarding_unit.reg_write_mem
+ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput101 net101 VGND VGND VPWR VPWR instruction_debug[23] sky130_fd_sc_hd__buf_8
Xoutput123 net123 VGND VGND VPWR VPWR pc_current[28] sky130_fd_sc_hd__buf_8
Xoutput112 net112 VGND VGND VPWR VPWR pc_current[17] sky130_fd_sc_hd__buf_8
Xoutput134 net134 VGND VGND VPWR VPWR pc_current[9] sky130_fd_sc_hd__buf_8
XFILLER_0_112_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1507_ _0496_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__clkbuf_4
X_1438_ net107 net415 _0458_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1369_ _0417_ _0419_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__or2b_1
XFILLER_0_37_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_90_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1223_ _0283_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_79_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1154_ _0780_ _0781_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__nand2_1
X_1085_ dmem.address\[12\] _0611_ _0613_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0938_ _0538_ net141 id_ex_rs2_data\[3\] VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_86 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0869_ _0524_ net335 VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1910_ clknet_leaf_1_clk net227 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dfxtp_2
X_1841_ clknet_leaf_2_clk _0157_ VGND VGND VPWR VPWR id_ex_rs2_data\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1772_ clknet_leaf_14_clk _0088_ VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1206_ _0829_ _0830_ _0564_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__a21oi_1
X_1137_ _0753_ _0765_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_101_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1068_ _0694_ _0700_ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_36_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_49_Left_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3 dmem.address\[7\] VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_58_Left_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1824_ clknet_leaf_9_clk _0140_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_13_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1755_ clknet_leaf_19_clk _0072_ VGND VGND VPWR VPWR forwarding_unit.rs2_ex\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1686_ clknet_leaf_20_clk _0003_ VGND VGND VPWR VPWR register_file.write_data\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_40_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1540_ net383 _0503_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1471_ _0564_ net461 _0482_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__nor3_1
XFILLER_0_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_Left_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_87_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1807_ clknet_leaf_9_clk net235 VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold211 net56 VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold200 id_alu_src\[0\] VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold233 _0099_ VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__dlygate4sd3_1
X_1738_ clknet_leaf_4_clk _0055_ VGND VGND VPWR VPWR dmem.address\[22\] sky130_fd_sc_hd__dfxtp_1
Xhold222 _0091_ VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold244 dmem.address\[13\] VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold266 _0481_ VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 _0100_ VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__dlygate4sd3_1
X_1669_ net337 _0592_ net535 VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__and3_1
Xhold277 _0439_ VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold299 register_file.write_data\[27\] VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 net1 VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0971_ register_file.write_data\[5\] id_ex_rs2_data\[5\] _0609_ VGND VGND VPWR VPWR
+ _0610_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1523_ net280 _0496_ _0498_ net83 VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1454_ net113 net463 _0468_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__and3_1
X_1385_ _0428_ _0434_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_124_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire1 net170 VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_53_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1170_ _0794_ _0795_ _0796_ _0613_ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_48_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0954_ _0568_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0885_ register_file.write_data\[0\] id_ex_rs1_data\[0\] _0528_ VGND VGND VPWR VPWR
+ _0529_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput124 net124 VGND VGND VPWR VPWR pc_current[29] sky130_fd_sc_hd__buf_8
XFILLER_0_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput113 net113 VGND VGND VPWR VPWR pc_current[18] sky130_fd_sc_hd__buf_8
Xoutput102 net102 VGND VGND VPWR VPWR instruction_debug[5] sky130_fd_sc_hd__buf_8
XFILLER_0_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput135 net135 VGND VGND VPWR VPWR pipeline_state[0] sky130_fd_sc_hd__buf_12
XFILLER_0_112_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1506_ net218 _0497_ _0499_ net388 VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__a22o_1
X_1437_ net457 _0458_ net415 VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__a21oi_1
X_1368_ net418 _0418_ _0692_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1299_ _0352_ _0354_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Left_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1222_ _0281_ _0282_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__or2_1
X_1153_ _0777_ _0779_ VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__or2_1
X_1084_ register_file.write_data\[12\] id_ex_rs2_data\[12\] _0609_ VGND VGND VPWR
+ VPWR _0716_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0937_ _0576_ _0577_ _0578_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_9_clk net177 VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0868_ _0524_ net370 VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1840_ clknet_leaf_2_clk _0156_ VGND VGND VPWR VPWR id_ex_rs2_data\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1771_ clknet_leaf_14_clk net504 VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1205_ _0819_ _0821_ _0817_ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1136_ _0594_ _0763_ _0764_ _0613_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1067_ _0694_ _0700_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold4 _0008_ VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1823_ clknet_leaf_9_clk _0139_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1754_ clknet_leaf_19_clk _0071_ VGND VGND VPWR VPWR forwarding_unit.rs2_ex\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1685_ clknet_leaf_20_clk _0002_ VGND VGND VPWR VPWR register_file.write_data\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_40_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_Right_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_127_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1119_ register_file.write_data\[14\] id_ex_rs2_data\[14\] _0609_ VGND VGND VPWR
+ VPWR _0749_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_4_Left_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1470_ net541 net460 _0478_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1806_ clknet_leaf_8_clk net247 VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold201 _0597_ VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold234 dmem.address\[31\] VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 dmem.address\[30\] VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 net57 VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__dlygate4sd3_1
X_1737_ clknet_leaf_4_clk _0054_ VGND VGND VPWR VPWR dmem.address\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold267 _0102_ VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 net93 VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 net112 VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold278 _0440_ VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1668_ net337 _0592_ net16 VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__and3_1
Xhold289 net124 VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1599_ net341 net314 _0507_ net343 VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0970_ _0566_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_43_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1522_ net278 _0496_ _0498_ net82 VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1453_ net113 _0468_ net463 VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1384_ _0431_ _0433_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_124_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire2 net171 VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__buf_1
XFILLER_0_111_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_85_Left_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_94_Left_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0953_ net522 _0591_ _0593_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0884_ _0527_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput114 net114 VGND VGND VPWR VPWR pc_current[19] sky130_fd_sc_hd__buf_8
Xoutput103 net103 VGND VGND VPWR VPWR instruction_debug[7] sky130_fd_sc_hd__buf_8
XFILLER_0_2_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput125 net125 VGND VGND VPWR VPWR pc_current[2] sky130_fd_sc_hd__buf_8
XFILLER_0_23_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput136 net136 VGND VGND VPWR VPWR pipeline_state[1] sky130_fd_sc_hd__buf_8
X_1505_ net210 _0497_ _0499_ net387 VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1436_ net457 _0458_ _0460_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__o21a_1
X_1367_ register_file.write_data\[30\] id_ex_rs1_data\[30\] _0690_ VGND VGND VPWR
+ VPWR _0418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1298_ net421 _0353_ _0692_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_48 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1221_ _0839_ _0840_ _0280_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1152_ _0777_ _0779_ VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1083_ _0713_ _0714_ _0715_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0936_ _0576_ _0577_ _0564_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0867_ _0524_ net380 VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1419_ net500 _0446_ _0449_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_3_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_129_Right_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XCPU_core_160 VGND VGND VPWR VPWR CPU_core_160/HI instruction_debug[28] sky130_fd_sc_hd__conb_1
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1770_ clknet_leaf_14_clk _0086_ VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1204_ _0826_ _0828_ VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__xnor2_2
X_1135_ dmem.address\[15\] _0611_ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1066_ _0697_ _0699_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0919_ _0553_ _0554_ _0560_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__nand3_1
XFILLER_0_16_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1899_ clknet_leaf_0_clk net211 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_70_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold5 dmem.address\[27\] VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_89_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1822_ clknet_leaf_9_clk net342 VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1753_ clknet_leaf_20_clk _0070_ VGND VGND VPWR VPWR forwarding_unit.rs1_ex\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1684_ clknet_leaf_20_clk _0001_ VGND VGND VPWR VPWR register_file.write_data\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_13_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1118_ _0747_ _0748_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1049_ _0664_ _0676_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_105_Left_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_74 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_114_Left_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1805_ clknet_leaf_9_clk net241 VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dfxtp_1
X_1736_ clknet_leaf_4_clk _0053_ VGND VGND VPWR VPWR dmem.address\[20\] sky130_fd_sc_hd__dfxtp_1
Xhold202 _0598_ VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold235 dmem.address\[24\] VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 net100 VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold224 net55 VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold268 net114 VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 _0094_ VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 forwarding_unit.rs2_ex\[1\] VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__dlygate4sd3_1
X_1667_ _0517_ _0518_ net524 VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_123_Left_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold279 net123 VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1598_ net351 net314 _0507_ net357 VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_132_Left_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1521_ net282 _0496_ _0498_ net81 VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1452_ net516 _0468_ _0470_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1383_ net429 _0432_ _0692_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_124_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1719_ clknet_leaf_20_clk net523 VGND VGND VPWR VPWR dmem.address\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire3 net172 VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__buf_1
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0952_ net522 _0591_ _0592_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0883_ net308 _0526_ forwarding_unit.rs1_ex\[0\] VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__or3b_1
XFILLER_0_125_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput115 net115 VGND VGND VPWR VPWR pc_current[20] sky130_fd_sc_hd__buf_8
XFILLER_0_11_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput104 net104 VGND VGND VPWR VPWR instruction_debug[8] sky130_fd_sc_hd__buf_8
XFILLER_0_2_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput126 net126 VGND VGND VPWR VPWR pc_current[30] sky130_fd_sc_hd__buf_8
Xoutput137 net137 VGND VGND VPWR VPWR pipeline_state[2] sky130_fd_sc_hd__buf_8
XFILLER_0_100_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1504_ net302 _0497_ _0499_ net394 VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1435_ net457 _0458_ _0564_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1366_ _0413_ _0416_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__xor2_1
XFILLER_0_128_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1297_ register_file.write_data\[25\] id_ex_rs1_data\[25\] _0690_ VGND VGND VPWR
+ VPWR _0353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1220_ _0839_ _0840_ _0280_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__a21oi_1
X_1151_ net376 _0778_ _0620_ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1082_ _0713_ _0714_ _0521_ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0935_ _0546_ net527 _0561_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0866_ _0524_ net374 VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_132_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1418_ net500 _0446_ _0564_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_3_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1349_ _0350_ _0365_ _0377_ _0390_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XCPU_core_150 VGND VGND VPWR VPWR CPU_core_150/HI instruction_debug[13] sky130_fd_sc_hd__conb_1
XCPU_core_161 VGND VGND VPWR VPWR CPU_core_161/HI instruction_debug[29] sky130_fd_sc_hd__conb_1
XFILLER_0_88_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1203_ net370 _0827_ _0692_ VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1134_ register_file.write_data\[15\] id_ex_rs2_data\[15\] _0609_ VGND VGND VPWR
+ VPWR _0763_ sky130_fd_sc_hd__mux2_1
X_1065_ _0658_ _0698_ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_101_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1898_ clknet_leaf_21_clk _0214_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dfxtp_1
X_0918_ _0553_ _0554_ net531 VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0849_ _0522_ _0523_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_8_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold6 _0028_ VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_27_Left_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1821_ clknet_leaf_9_clk net352 VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_10_clk net178 VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_8
X_1752_ clknet_leaf_16_clk _0069_ VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_13_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1683_ _0440_ _0443_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_36_Left_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_84 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1117_ _0725_ _0734_ _0746_ _0607_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__a31o_1
X_1048_ _0681_ _0682_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_560 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_clk net174 VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1804_ clknet_leaf_7_clk _0120_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_74 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1735_ clknet_leaf_4_clk _0052_ VGND VGND VPWR VPWR dmem.address\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold214 net19 VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold203 _0601_ VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 dmem.address\[10\] VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 if_id_valid VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 net92 VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 _0471_ VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 net65 VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1666_ _0517_ _0518_ net14 VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__and3_1
X_1597_ net494 net314 _0507_ net347 VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1520_ net222 _0500_ _0501_ net250 VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1451_ net516 _0468_ _0564_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__a21oi_1
X_1382_ register_file.write_data\[31\] id_ex_rs1_data\[31\] _0690_ VGND VGND VPWR
+ VPWR _0432_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1718_ clknet_leaf_20_clk net532 VGND VGND VPWR VPWR dmem.address\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1649_ _0441_ _0411_ net260 VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__and3_1
Xwire4 clk VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0951_ _0519_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__buf_1
XFILLER_0_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0882_ net313 net308 net386 VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput116 net116 VGND VGND VPWR VPWR pc_current[21] sky130_fd_sc_hd__buf_8
XFILLER_0_11_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput105 net105 VGND VGND VPWR VPWR pc_current[10] sky130_fd_sc_hd__buf_8
XFILLER_0_51_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput127 net127 VGND VGND VPWR VPWR pc_current[31] sky130_fd_sc_hd__buf_8
XFILLER_0_121_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput138 net138 VGND VGND VPWR VPWR pipeline_state[3] sky130_fd_sc_hd__buf_8
X_1503_ net296 _0497_ _0499_ net391 VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__a22o_1
X_1434_ net498 _0457_ _0459_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_52_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1365_ _0837_ _0415_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1296_ _0350_ _0351_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1150_ register_file.write_data\[16\] id_ex_rs1_data\[16\] _0618_ VGND VGND VPWR
+ VPWR _0778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1081_ _0689_ _0693_ _0702_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_99_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0934_ _0573_ _0575_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0865_ _0524_ net376 VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1417_ _0446_ _0448_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1348_ _0391_ _0393_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_3_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1279_ register_file.write_data\[24\] id_ex_rs2_data\[24\] _0833_ VGND VGND VPWR
+ VPWR _0336_ sky130_fd_sc_hd__mux2_1
Xwire20 clknet_1_1__leaf_clk VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_78_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XCPU_core_151 VGND VGND VPWR VPWR CPU_core_151/HI instruction_debug[14] sky130_fd_sc_hd__conb_1
XCPU_core_162 VGND VGND VPWR VPWR CPU_core_162/HI instruction_debug[30] sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_110_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1202_ register_file.write_data\[19\] id_ex_rs1_data\[19\] _0690_ VGND VGND VPWR
+ VPWR _0827_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1133_ _0754_ _0756_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__or2b_1
X_1064_ _0668_ _0680_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0917_ _0523_ _0556_ _0557_ _0559_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1897_ clknet_leaf_21_clk _0213_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0848_ net411 VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold7 register_file.write_data\[19\] VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1820_ clknet_leaf_9_clk net470 VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1751_ clknet_leaf_19_clk _0068_ VGND VGND VPWR VPWR forwarding_unit.rd_wb\[1\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_52_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1682_ net330 _0275_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__nor2b_1
XFILLER_0_53_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_127_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1116_ _0725_ _0734_ _0746_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1047_ _0671_ _0670_ _0680_ _0607_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__a31o_1
XFILLER_0_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_122_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1949_ clknet_leaf_5_clk _0265_ VGND VGND VPWR VPWR id_ex_rs1_data\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1803_ clknet_leaf_7_clk _0119_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1734_ clknet_leaf_4_clk _0051_ VGND VGND VPWR VPWR dmem.address\[18\] sky130_fd_sc_hd__dfxtp_1
Xhold215 register_file.write_data\[26\] VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 dmem.address\[25\] VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 _0626_ VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold248 net90 VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 net91 VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold237 dmem.address\[5\] VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__dlygate4sd3_1
X_1665_ _0517_ _0518_ net364 VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__and3_1
X_1596_ net280 net314 _0507_ net349 VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_55_Left_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Left_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1450_ net451 _0467_ _0469_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1381_ _0794_ _0429_ _0430_ _0837_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_124_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1717_ clknet_leaf_20_clk net529 VGND VGND VPWR VPWR ex_mem_alu_result\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1648_ _0441_ _0411_ net264 VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire5 clknet_0_clk VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__buf_1
X_1579_ net218 _0506_ _0508_ net276 VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_68_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_72_Left_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0950_ _0576_ _0577_ _0590_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0881_ _0525_ net429 VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_124_Right_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_81_Left_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput106 net106 VGND VGND VPWR VPWR pc_current[11] sky130_fd_sc_hd__buf_8
Xoutput117 net117 VGND VGND VPWR VPWR pc_current[22] sky130_fd_sc_hd__buf_8
X_1502_ register_file.write_data\[7\] _0497_ _0499_ net446 VGND VGND VPWR VPWR _0116_
+ sky130_fd_sc_hd__a22o_1
Xoutput128 net128 VGND VGND VPWR VPWR pc_current[3] sky130_fd_sc_hd__buf_8
XFILLER_0_23_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1433_ _0452_ _0458_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_52_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1364_ net418 _0414_ _0835_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1295_ _0317_ _0320_ _0338_ _0348_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__o31ai_1
XPHY_EDGE_ROW_90_Left_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_129_Left_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1080_ _0711_ _0712_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0933_ net422 _0574_ _0532_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0864_ _0524_ net385 VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_132_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1416_ _0592_ net402 VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__nand2_1
X_1347_ _0394_ _0397_ _0399_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_3_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire10 net182 VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__buf_1
XFILLER_0_78_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1278_ _0317_ _0320_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire21 net195 VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__buf_1
XFILLER_0_78_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XCPU_core_152 VGND VGND VPWR VPWR CPU_core_152/HI instruction_debug[16] sky130_fd_sc_hd__conb_1
XCPU_core_163 VGND VGND VPWR VPWR CPU_core_163/HI instruction_debug[31] sky130_fd_sc_hd__conb_1
XFILLER_0_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1201_ _0813_ _0825_ VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__xor2_2
X_1132_ _0628_ _0760_ _0761_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__and3_1
X_1063_ _0671_ _0695_ _0696_ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0916_ register_file.write_data\[1\] _0558_ _0556_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_116_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1896_ clknet_leaf_21_clk _0212_ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0847_ _0521_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__buf_1
XFILLER_0_70_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold8 _0224_ VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1750_ clknet_leaf_19_clk _0067_ VGND VGND VPWR VPWR forwarding_unit.rd_wb\[0\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_4_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1681_ _0443_ _0275_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__nor2b_1
XFILLER_0_13_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1115_ _0744_ _0745_ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__or2b_1
XFILLER_0_45_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1046_ _0671_ _0670_ _0680_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1948_ clknet_leaf_5_clk _0264_ VGND VGND VPWR VPWR id_ex_rs1_data\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1879_ clknet_leaf_6_clk net305 VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1802_ clknet_leaf_7_clk _0118_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1733_ clknet_leaf_4_clk _0050_ VGND VGND VPWR VPWR dmem.address\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold216 ex_mem_alu_result\[1\] VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__dlygate4sd3_1
Xhold205 _0038_ VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 net76 VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 dmem.address\[2\] VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold238 forwarding_unit.reg_write_mem VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__dlygate4sd3_1
X_1664_ _0517_ _0518_ net519 VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__and3_1
X_1595_ net278 net314 _0507_ net50 VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1029_ _0660_ _0664_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_101_Left_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_110_Left_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1380_ net429 _0835_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_124_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1716_ clknet_leaf_20_clk net509 VGND VGND VPWR VPWR ex_mem_alu_result\[0\] sky130_fd_sc_hd__dfxtp_1
X_1647_ _0441_ _0411_ net477 VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire6 _0536_ VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__buf_1
X_1578_ net210 _0506_ _0508_ net270 VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0880_ _0525_ net418 VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput107 net107 VGND VGND VPWR VPWR pc_current[12] sky130_fd_sc_hd__buf_8
Xoutput118 net118 VGND VGND VPWR VPWR pc_current[23] sky130_fd_sc_hd__buf_8
X_1501_ register_file.write_data\[6\] _0497_ _0499_ net440 VGND VGND VPWR VPWR _0115_
+ sky130_fd_sc_hd__a22o_1
Xoutput129 net129 VGND VGND VPWR VPWR pc_current[4] sky130_fd_sc_hd__buf_8
XFILLER_0_50_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1432_ net502 net505 net498 _0453_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_52_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1363_ register_file.write_data\[30\] id_ex_rs2_data\[30\] _0833_ VGND VGND VPWR
+ VPWR _0414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1294_ _0349_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_108_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_22 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0932_ register_file.write_data\[2\] id_ex_rs1_data\[2\] _0528_ VGND VGND VPWR VPWR
+ _0574_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0863_ _0524_ net382 VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1415_ net129 net330 net125 net401 VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__a31o_1
XFILLER_0_48_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1346_ _0521_ _0398_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_3_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1277_ _0313_ _0330_ _0331_ _0288_ _0333_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__a221oi_2
Xwire11 net180 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__dlymetal6s2s_1
Xwire22 net191 VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__buf_1
XFILLER_0_78_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XCPU_core_153 VGND VGND VPWR VPWR CPU_core_153/HI instruction_debug[17] sky130_fd_sc_hd__conb_1
XFILLER_0_15_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XCPU_core_164 VGND VGND VPWR VPWR CPU_core_164/HI pc_current[0] sky130_fd_sc_hd__conb_1
XFILLER_0_30_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1200_ _0794_ _0823_ _0824_ _0613_ VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__o211a_1
X_1131_ _0757_ _0759_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__or2_1
X_1062_ _0677_ _0679_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_13_clk net191 VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_60_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0915_ forwarding_unit.rd_wb\[1\] _0538_ forwarding_unit.rs1_ex\[0\] VGND VGND VPWR
+ VPWR _0558_ sky130_fd_sc_hd__and3b_2
XFILLER_0_114_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1895_ clknet_leaf_21_clk _0211_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_116_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0846_ reset VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__buf_1
XFILLER_0_101_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1329_ _0378_ _0379_ _0382_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold9 register_file.write_data\[15\] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_89_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1680_ net434 net473 VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap139 _0623_ VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_2_clk net180 VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_119_Right_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1114_ _0739_ _0740_ _0743_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1045_ _0677_ _0679_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1947_ clknet_leaf_5_clk _0263_ VGND VGND VPWR VPWR id_ex_rs1_data\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1878_ clknet_leaf_6_clk net317 VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1801_ clknet_leaf_7_clk _0117_ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1732_ clknet_leaf_4_clk _0049_ VGND VGND VPWR VPWR dmem.address\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold217 ex_mem_valid VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold206 net130 VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__dlygate4sd3_1
X_1663_ _0517_ _0518_ net10 VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold239 net125 VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 dmem.address\[8\] VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__dlygate4sd3_1
X_1594_ net282 net314 _0507_ net318 VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1028_ _0568_ _0661_ _0662_ _0663_ _0543_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__o311a_1
XFILLER_0_48_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1715_ clknet_leaf_10_clk _0032_ VGND VGND VPWR VPWR register_file.write_data\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1646_ _0441_ _0411_ net486 VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire7 net176 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__dlymetal6s2s_1
X_1577_ net302 _0506_ _0508_ net64 VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput119 net119 VGND VGND VPWR VPWR pc_current[24] sky130_fd_sc_hd__buf_8
X_1500_ register_file.write_data\[5\] _0497_ _0499_ net453 VGND VGND VPWR VPWR _0114_
+ sky130_fd_sc_hd__a22o_1
Xoutput108 net108 VGND VGND VPWR VPWR pc_current[13] sky130_fd_sc_hd__buf_8
XFILLER_0_11_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1431_ _0522_ net503 _0457_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__nor3_1
XFILLER_0_120_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1362_ _0401_ _0404_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__nor2_1
Xoutput90 net90 VGND VGND VPWR VPWR debug_reg3[3] sky130_fd_sc_hd__buf_8
X_1293_ _0317_ _0320_ _0338_ _0348_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__or4_1
XFILLER_0_37_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_108_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1629_ net226 _0515_ _0516_ net14 VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0931_ _0553_ _0572_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__xor2_1
XFILLER_0_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0862_ _0524_ net439 VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_132_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1414_ net525 net401 net330 net125 VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__and4_1
XFILLER_0_48_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1345_ _0394_ _0397_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1276_ _0321_ _0323_ _0332_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_65_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire23 net193 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XCPU_core_143 VGND VGND VPWR VPWR CPU_core_143/HI instruction_debug[2] sky130_fd_sc_hd__conb_1
XCPU_core_154 VGND VGND VPWR VPWR CPU_core_154/HI instruction_debug[18] sky130_fd_sc_hd__conb_1
XFILLER_0_30_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XCPU_core_165 VGND VGND VPWR VPWR CPU_core_165/HI pc_current[1] sky130_fd_sc_hd__conb_1
XFILLER_0_100_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1130_ _0757_ _0759_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_129_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1061_ _0677_ _0679_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Left_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0914_ net530 _0528_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__nand2_1
X_1894_ clknet_leaf_21_clk _0210_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0845_ net424 _0520_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_116_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_87_Left_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1328_ _0381_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__inv_2
X_1259_ _0773_ _0832_ _0306_ _0294_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__or4b_2
XFILLER_0_39_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_96_Left_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1113_ _0739_ _0740_ _0743_ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1044_ net425 _0678_ _0620_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1946_ clknet_leaf_6_clk _0262_ VGND VGND VPWR VPWR id_ex_rs1_data\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1877_ clknet_leaf_6_clk net321 VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1800_ clknet_leaf_7_clk _0116_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1731_ clknet_leaf_4_clk _0048_ VGND VGND VPWR VPWR dmem.address\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold207 _0447_ VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__dlygate4sd3_1
X_1662_ _0517_ _0518_ net363 VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold218 id_ex_valid VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 ex_mem_alu_result\[0\] VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__dlygate4sd3_1
X_1593_ net222 _0509_ _0510_ net306 VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1027_ dmem.address\[8\] _0530_ _0567_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__or3_1
XFILLER_0_48_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1929_ clknet_leaf_0_clk net265 VGND VGND VPWR VPWR id_ex_rs1_data\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Left_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_24_Left_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Left_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Left_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold90 _0248_ VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_55 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_51_Left_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1714_ clknet_leaf_10_clk _0031_ VGND VGND VPWR VPWR register_file.write_data\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1645_ _0441_ _0411_ net501 VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1576_ net296 _0506_ _0508_ net63 VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__a22o_1
Xwire8 net184 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_60_Left_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput109 net109 VGND VGND VPWR VPWR pc_current[14] sky130_fd_sc_hd__buf_8
XFILLER_0_11_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput1 net1 VGND VGND VPWR VPWR debug_reg1[0] sky130_fd_sc_hd__buf_8
X_1430_ net502 net505 _0453_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1361_ _0405_ _0407_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_52_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput80 net80 VGND VGND VPWR VPWR debug_reg3[23] sky130_fd_sc_hd__buf_8
Xoutput91 net91 VGND VGND VPWR VPWR debug_reg3[4] sky130_fd_sc_hd__buf_8
X_1292_ _0794_ _0346_ _0347_ _0837_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_108_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1628_ net228 _0515_ _0516_ net13 VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__a22o_1
X_1559_ net347 net140 VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_107_Left_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_116_Left_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0930_ _0543_ _0570_ _0571_ _0534_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__a31o_1
XFILLER_0_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0861_ _0519_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__buf_1
XFILLER_0_36_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1413_ net331 _0445_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1344_ _0360_ _0362_ _0395_ _0396_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__a31o_1
X_1275_ _0307_ _0309_ _0321_ _0323_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__a22o_1
Xwire13 net182 VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__buf_1
XFILLER_0_64_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XCPU_core_144 VGND VGND VPWR VPWR CPU_core_144/HI instruction_debug[3] sky130_fd_sc_hd__conb_1
XFILLER_0_15_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XCPU_core_166 VGND VGND VPWR VPWR instruction_debug[0] CPU_core_166/LO sky130_fd_sc_hd__conb_1
XCPU_core_155 VGND VGND VPWR VPWR CPU_core_155/HI instruction_debug[19] sky130_fd_sc_hd__conb_1
XFILLER_0_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1060_ _0689_ _0693_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__xor2_2
XFILLER_0_88_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1962_ clknet_leaf_16_clk _0278_ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_28_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0913_ _0555_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__buf_2
X_1893_ clknet_leaf_21_clk _0209_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0844_ _0519_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__buf_1
XFILLER_0_43_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1327_ net200 _0380_ _0692_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__mux2_1
X_1258_ _0628_ _0315_ _0316_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__and3_1
X_1189_ register_file.write_data\[18\] id_ex_rs1_data\[18\] _0618_ VGND VGND VPWR
+ VPWR _0815_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_133_Right_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_111_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1112_ net439 _0556_ _0742_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__a21oi_1
X_1043_ register_file.write_data\[9\] id_ex_rs1_data\[9\] _0618_ VGND VGND VPWR VPWR
+ _0678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1945_ clknet_leaf_3_clk _0261_ VGND VGND VPWR VPWR id_ex_rs1_data\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1876_ clknet_leaf_6_clk net253 VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1730_ clknet_leaf_4_clk _0047_ VGND VGND VPWR VPWR dmem.address\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold208 _0082_ VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__dlygate4sd3_1
X_1661_ _0517_ _0518_ net8 VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__and3_1
Xhold219 dmem.address\[11\] VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1592_ net224 _0509_ _0510_ net304 VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1026_ _0526_ _0541_ id_ex_rs2_data\[8\] VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1928_ clknet_leaf_21_clk _0244_ VGND VGND VPWR VPWR id_ex_rs1_data\[4\] sky130_fd_sc_hd__dfxtp_1
X_1859_ clknet_leaf_1_clk net291 VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_40_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold91 net78 VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 _0186_ VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1713_ clknet_leaf_10_clk _0030_ VGND VGND VPWR VPWR register_file.write_data\[29\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_130_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1644_ _0441_ _0411_ net478 VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1575_ net481 _0506_ _0508_ net368 VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__a22o_1
Xwire9 net178 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_83_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1009_ _0584_ _0615_ _0645_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__nor3_2
XFILLER_0_76_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput2 net2 VGND VGND VPWR VPWR debug_reg1[10] sky130_fd_sc_hd__buf_12
XFILLER_0_120_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput70 net70 VGND VGND VPWR VPWR debug_reg3[14] sky130_fd_sc_hd__buf_8
X_1360_ _0519_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_52_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput81 net81 VGND VGND VPWR VPWR debug_reg3[24] sky130_fd_sc_hd__buf_8
Xoutput92 net92 VGND VGND VPWR VPWR debug_reg3[5] sky130_fd_sc_hd__buf_8
X_1291_ dmem.address\[25\] _0835_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_108_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1627_ net202 _0515_ _0516_ net11 VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1558_ net349 net140 VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__and2_1
X_1489_ _0493_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0860_ _0000_ net438 VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1412_ net129 net330 net125 _0521_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_114_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1343_ _0370_ _0384_ _0383_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__a21oi_1
X_1274_ _0284_ _0301_ _0327_ _0324_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__nor4_1
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire25 net194 VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_16_clk net189 VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_19_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0989_ net399 _0627_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XCPU_core_145 VGND VGND VPWR VPWR CPU_core_145/HI instruction_debug[6] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_76_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XCPU_core_167 VGND VGND VPWR VPWR instruction_debug[1] CPU_core_167/LO sky130_fd_sc_hd__conb_1
XCPU_core_156 VGND VGND VPWR VPWR CPU_core_156/HI instruction_debug[24] sky130_fd_sc_hd__conb_1
XFILLER_0_30_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_114_Right_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1961_ clknet_leaf_16_clk _0277_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1892_ clknet_leaf_21_clk _0208_ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dfxtp_1
X_0912_ forwarding_unit.rd_mem\[1\] forwarding_unit.rs1_ex\[0\] _0535_ VGND VGND VPWR
+ VPWR _0555_ sky130_fd_sc_hd__and3b_1
XFILLER_0_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0843_ _0519_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__buf_1
XFILLER_0_43_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_5_clk net182 VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_58_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1326_ register_file.write_data\[27\] id_ex_rs1_data\[27\] _0690_ VGND VGND VPWR
+ VPWR _0380_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1257_ _0313_ _0314_ _0312_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1188_ _0793_ _0798_ _0811_ VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_111_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1111_ id_ex_rs1_data\[13\] _0558_ _0741_ _0532_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap1 _0539_ VGND VGND VPWR VPWR net542 sky130_fd_sc_hd__clkbuf_1
X_1042_ _0672_ _0676_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_122_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1944_ clknet_leaf_0_clk _0260_ VGND VGND VPWR VPWR id_ex_rs1_data\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1875_ clknet_leaf_6_clk net267 VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1309_ net324 _0835_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire140 net405 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_4
X_1660_ _0517_ _0518_ net7 VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__and3_1
XFILLER_0_111_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1591_ net226 _0509_ _0510_ net316 VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__a22o_1
Xhold209 net101 VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1025_ register_file.write_data\[8\] _0538_ net542 VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1927_ clknet_leaf_21_clk _0243_ VGND VGND VPWR VPWR id_ex_rs1_data\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1858_ clknet_leaf_1_clk net295 VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_114_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1789_ clknet_leaf_12_clk net476 VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold92 _0130_ VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 net35 VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 _0245_ VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_133_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1712_ clknet_leaf_10_clk _0029_ VGND VGND VPWR VPWR register_file.write_data\[28\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_81_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1643_ _0441_ _0411_ net483 VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1574_ net482 _0506_ _0508_ net366 VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1008_ _0631_ _0644_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_81_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_128_Right_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput3 net3 VGND VGND VPWR VPWR debug_reg1[11] sky130_fd_sc_hd__buf_12
XFILLER_0_50_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput60 net60 VGND VGND VPWR VPWR debug_reg2[5] sky130_fd_sc_hd__buf_8
XFILLER_0_128_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput82 net82 VGND VGND VPWR VPWR debug_reg3[25] sky130_fd_sc_hd__buf_8
Xoutput71 net71 VGND VGND VPWR VPWR debug_reg3[15] sky130_fd_sc_hd__buf_8
Xoutput93 net93 VGND VGND VPWR VPWR debug_reg3[6] sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_52_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1290_ register_file.write_data\[25\] id_ex_rs2_data\[25\] _0833_ VGND VGND VPWR
+ VPWR _0346_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1626_ net216 _0515_ _0516_ net10 VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1557_ net539 net140 VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1488_ _0526_ reset mem_wb_valid VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__or3b_4
XFILLER_0_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1411_ net330 net125 net129 VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_39_Left_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1342_ _0369_ _0384_ _0383_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__a21oi_1
X_1273_ _0327_ _0324_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire15 clknet_1_0__leaf_clk VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_48_Left_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0988_ net398 _0606_ _0625_ _0607_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__a31o_1
XFILLER_0_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_57_Left_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XCPU_core_146 VGND VGND VPWR VPWR CPU_core_146/HI instruction_debug[9] sky130_fd_sc_hd__conb_1
XCPU_core_168 VGND VGND VPWR VPWR instruction_debug[4] CPU_core_168/LO sky130_fd_sc_hd__conb_1
XCPU_core_157 VGND VGND VPWR VPWR CPU_core_157/HI instruction_debug[25] sky130_fd_sc_hd__conb_1
XFILLER_0_30_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1609_ net292 _0512_ _0514_ net486 VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1960_ clknet_leaf_18_clk _0276_ VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_55_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1891_ clknet_leaf_21_clk _0207_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dfxtp_1
X_0911_ _0534_ _0544_ _0548_ _0552_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_50_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0842_ reset VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1325_ _0350_ _0365_ _0377_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_71_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1256_ _0312_ _0313_ _0314_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__or3_1
XFILLER_0_78_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1187_ _0773_ _0812_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1110_ register_file.write_data\[13\] _0528_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1041_ _0568_ _0673_ _0674_ _0675_ _0543_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__o311a_1
XFILLER_0_88_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_122_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1943_ clknet_leaf_2_clk _0259_ VGND VGND VPWR VPWR id_ex_rs1_data\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1874_ clknet_leaf_6_clk net269 VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1308_ register_file.write_data\[26\] id_ex_rs2_data\[26\] _0833_ VGND VGND VPWR
+ VPWR _0363_ sky130_fd_sc_hd__mux2_1
X_1239_ _0295_ _0296_ _0298_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_84_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1590_ net228 _0509_ _0510_ net320 VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1024_ _0659_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__buf_2
XFILLER_0_49_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1926_ clknet_leaf_20_clk _0242_ VGND VGND VPWR VPWR id_ex_rs1_data\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1857_ clknet_leaf_1_clk net301 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_114_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1788_ clknet_leaf_12_clk _0104_ VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_109_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold71 net42 VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 _0189_ VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 _0184_ VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 net77 VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_11_Left_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1711_ clknet_leaf_8_clk net201 VGND VGND VPWR VPWR register_file.write_data\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1642_ net337 _0521_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_20_Left_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1573_ register_file.write_data\[5\] _0506_ _0508_ net488 VGND VGND VPWR VPWR _0178_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1007_ _0594_ _0642_ _0643_ _0543_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1909_ clknet_leaf_1_clk net229 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_130_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput4 net4 VGND VGND VPWR VPWR debug_reg1[12] sky130_fd_sc_hd__buf_12
XFILLER_0_120_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput50 net50 VGND VGND VPWR VPWR debug_reg2[25] sky130_fd_sc_hd__buf_8
Xoutput61 net61 VGND VGND VPWR VPWR debug_reg2[6] sky130_fd_sc_hd__buf_8
XFILLER_0_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput83 net83 VGND VGND VPWR VPWR debug_reg3[26] sky130_fd_sc_hd__buf_8
XFILLER_0_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput72 net72 VGND VGND VPWR VPWR debug_reg3[16] sky130_fd_sc_hd__buf_8
Xoutput94 net94 VGND VGND VPWR VPWR debug_reg3[7] sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_52_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1625_ net214 _0515_ _0516_ net9 VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__a22o_1
X_1556_ net318 net140 VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1487_ net497 _0490_ _0492_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_418 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1410_ _0522_ _0443_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1341_ _0391_ _0393_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__xnor2_1
X_1272_ _0784_ _0789_ _0285_ _0328_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__a211o_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_55 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0987_ net398 _0606_ _0625_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_131_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XCPU_core_147 VGND VGND VPWR VPWR CPU_core_147/HI instruction_debug[10] sky130_fd_sc_hd__conb_1
XCPU_core_158 VGND VGND VPWR VPWR CPU_core_158/HI instruction_debug[26] sky130_fd_sc_hd__conb_1
XFILLER_0_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1608_ net290 _0512_ _0514_ net501 VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1539_ net537 _0503_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold190 dmem.address\[15\] VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0910_ _0548_ _0552_ _0534_ _0544_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__a211o_1
XFILLER_0_126_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1890_ clknet_leaf_21_clk _0206_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1324_ _0350_ _0365_ _0377_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__or3_1
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1255_ _0284_ _0289_ _0301_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__nor3_1
XPHY_EDGE_ROW_3_Left_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1186_ _0798_ _0811_ VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1040_ dmem.address\[9\] _0530_ _0567_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__or3_1
XFILLER_0_88_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1942_ clknet_leaf_3_clk _0258_ VGND VGND VPWR VPWR id_ex_rs1_data\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1873_ clknet_leaf_6_clk net255 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_12_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1307_ _0355_ _0361_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__nor2_1
X_1238_ net322 _0297_ _0620_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1169_ dmem.address\[17\] _0611_ VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_590 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_Left_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_84_Left_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1023_ _0584_ _0615_ _0645_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_93_Left_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1925_ clknet_leaf_21_clk _0241_ VGND VGND VPWR VPWR id_ex_rs1_data\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1856_ clknet_leaf_8_clk _0172_ VGND VGND VPWR VPWR id_ex_rs2_data\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1787_ clknet_leaf_12_clk net456 VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold50 _0127_ VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 register_file.write_data\[25\] VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 _0191_ VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 net39 VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold94 _0129_ VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1710_ clknet_leaf_5_clk net325 VGND VGND VPWR VPWR register_file.write_data\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1641_ _0522_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1572_ register_file.write_data\[4\] _0506_ _0508_ net389 VGND VGND VPWR VPWR _0177_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1006_ dmem.address\[7\] _0537_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_81_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1908_ clknet_leaf_1_clk net203 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_115_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1839_ clknet_leaf_2_clk _0155_ VGND VGND VPWR VPWR id_ex_rs2_data\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_20_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput5 net5 VGND VGND VPWR VPWR debug_reg1[13] sky130_fd_sc_hd__buf_12
Xoutput51 net51 VGND VGND VPWR VPWR debug_reg2[26] sky130_fd_sc_hd__buf_8
Xoutput40 net40 VGND VGND VPWR VPWR debug_reg2[16] sky130_fd_sc_hd__buf_8
XFILLER_0_120_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput84 net84 VGND VGND VPWR VPWR debug_reg3[27] sky130_fd_sc_hd__buf_8
Xoutput73 net73 VGND VGND VPWR VPWR debug_reg3[17] sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_52_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput62 net62 VGND VGND VPWR VPWR debug_reg2[7] sky130_fd_sc_hd__buf_8
Xoutput95 net95 VGND VGND VPWR VPWR debug_reg3[8] sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_8_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1624_ net206 _0515_ _0516_ net8 VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1555_ net306 _0504_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__and2_1
X_1486_ net497 _0490_ _0452_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_19_clk net176 VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1340_ net435 _0392_ _0692_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__mux2_1
X_1271_ _0284_ _0301_ _0327_ _0324_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire17 net187 VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__buf_1
XFILLER_0_74_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0986_ _0622_ _0624_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_8_clk net177 VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_76_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XCPU_core_148 VGND VGND VPWR VPWR CPU_core_148/HI instruction_debug[11] sky130_fd_sc_hd__conb_1
XCPU_core_159 VGND VGND VPWR VPWR CPU_core_159/HI instruction_debug[27] sky130_fd_sc_hd__conb_1
X_1607_ net294 _0512_ _0514_ net478 VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1538_ net368 _0503_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1469_ net119 _0478_ net460 VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_2_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold180 _0018_ VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold191 forwarding_unit.reg_write_wb VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1323_ _0376_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_71_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1254_ _0281_ _0300_ _0299_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__a21o_1
X_1185_ _0613_ _0810_ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_104_Left_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0969_ _0606_ _0608_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_113_Left_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_122_Left_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_131_Left_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1941_ clknet_leaf_0_clk _0257_ VGND VGND VPWR VPWR id_ex_rs1_data\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1872_ clknet_leaf_6_clk net257 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1306_ _0345_ _0356_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__and2b_1
XFILLER_0_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1237_ register_file.write_data\[21\] id_ex_rs1_data\[21\] _0618_ VGND VGND VPWR
+ VPWR _0297_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1168_ register_file.write_data\[17\] id_ex_rs2_data\[17\] _0609_ VGND VGND VPWR
+ VPWR _0795_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_84_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1099_ _0694_ _0697_ _0712_ _0729_ _0730_ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__a311oi_2
XFILLER_0_75_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1022_ net139 _0637_ _0638_ _0653_ _0657_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__o41a_2
XFILLER_0_88_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1924_ clknet_leaf_20_clk _0240_ VGND VGND VPWR VPWR id_ex_rs1_data\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1855_ clknet_leaf_8_clk _0171_ VGND VGND VPWR VPWR id_ex_rs2_data\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1786_ clknet_leaf_12_clk net462 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_123_Right_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold40 _0123_ VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 net69 VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 net41 VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 _0188_ VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 _0134_ VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 register_file.write_data\[2\] VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_133_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1640_ _0442_ net510 VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1571_ net292 _0506_ _0508_ net58 VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1005_ register_file.write_data\[7\] id_ex_rs2_data\[7\] _0566_ VGND VGND VPWR VPWR
+ _0642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1907_ clknet_leaf_1_clk net217 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_45_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1838_ clknet_leaf_2_clk _0154_ VGND VGND VPWR VPWR id_ex_rs2_data\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1769_ clknet_leaf_14_clk net493 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput6 net6 VGND VGND VPWR VPWR debug_reg1[14] sky130_fd_sc_hd__buf_12
XFILLER_0_31_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput52 net52 VGND VGND VPWR VPWR debug_reg2[27] sky130_fd_sc_hd__buf_8
Xoutput41 net41 VGND VGND VPWR VPWR debug_reg2[17] sky130_fd_sc_hd__buf_8
Xoutput30 net30 VGND VGND VPWR VPWR debug_reg1[7] sky130_fd_sc_hd__buf_8
Xoutput85 net85 VGND VGND VPWR VPWR debug_reg3[28] sky130_fd_sc_hd__buf_8
Xoutput74 net74 VGND VGND VPWR VPWR debug_reg3[18] sky130_fd_sc_hd__buf_8
Xoutput63 net63 VGND VGND VPWR VPWR debug_reg2[8] sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_52_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput96 net96 VGND VGND VPWR VPWR debug_reg3[9] sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_8_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_26 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1623_ net204 _0515_ _0516_ net7 VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1554_ net304 _0504_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1485_ net479 _0488_ _0491_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__o21a_1
.ends

