module CPU_core (clk,
    reset,
    debug_reg1,
    debug_reg2,
    debug_reg3,
    instruction_debug,
    pc_current,
    pipeline_state);
 input clk;
 input reset;
 output [31:0] debug_reg1;
 output [31:0] debug_reg2;
 output [31:0] debug_reg3;
 output [31:0] instruction_debug;
 output [31:0] pc_current;
 output [3:0] pipeline_state;

 wire net166;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net167;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net143;
 wire net162;
 wire net163;
 wire net144;
 wire net168;
 wire net145;
 wire net146;
 wire net164;
 wire net165;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire \dmem.address[10] ;
 wire \dmem.address[11] ;
 wire \dmem.address[12] ;
 wire \dmem.address[13] ;
 wire \dmem.address[14] ;
 wire \dmem.address[15] ;
 wire \dmem.address[16] ;
 wire \dmem.address[17] ;
 wire \dmem.address[18] ;
 wire \dmem.address[19] ;
 wire \dmem.address[20] ;
 wire \dmem.address[21] ;
 wire \dmem.address[22] ;
 wire \dmem.address[23] ;
 wire \dmem.address[24] ;
 wire \dmem.address[25] ;
 wire \dmem.address[26] ;
 wire \dmem.address[27] ;
 wire \dmem.address[28] ;
 wire \dmem.address[29] ;
 wire \dmem.address[2] ;
 wire \dmem.address[30] ;
 wire \dmem.address[31] ;
 wire \dmem.address[3] ;
 wire \dmem.address[4] ;
 wire \dmem.address[5] ;
 wire \dmem.address[6] ;
 wire \dmem.address[7] ;
 wire \dmem.address[8] ;
 wire \dmem.address[9] ;
 wire \ex_mem_alu_result[0] ;
 wire \ex_mem_alu_result[1] ;
 wire ex_mem_valid;
 wire \forwarding_unit.rd_mem[0] ;
 wire \forwarding_unit.rd_mem[1] ;
 wire \forwarding_unit.rd_wb[0] ;
 wire \forwarding_unit.rd_wb[1] ;
 wire \forwarding_unit.reg_write_mem ;
 wire \forwarding_unit.reg_write_wb ;
 wire \forwarding_unit.rs1_ex[0] ;
 wire \forwarding_unit.rs2_ex[0] ;
 wire \forwarding_unit.rs2_ex[1] ;
 wire \forwarding_unit.rs2_ex[3] ;
 wire \id_alu_src[0] ;
 wire \id_ex_immediate[0] ;
 wire \id_ex_immediate[1] ;
 wire \id_ex_immediate[3] ;
 wire \id_ex_rd_addr[0] ;
 wire \id_ex_rs1_data[0] ;
 wire \id_ex_rs1_data[10] ;
 wire \id_ex_rs1_data[11] ;
 wire \id_ex_rs1_data[12] ;
 wire \id_ex_rs1_data[13] ;
 wire \id_ex_rs1_data[14] ;
 wire \id_ex_rs1_data[15] ;
 wire \id_ex_rs1_data[16] ;
 wire \id_ex_rs1_data[17] ;
 wire \id_ex_rs1_data[18] ;
 wire \id_ex_rs1_data[19] ;
 wire \id_ex_rs1_data[1] ;
 wire \id_ex_rs1_data[20] ;
 wire \id_ex_rs1_data[21] ;
 wire \id_ex_rs1_data[22] ;
 wire \id_ex_rs1_data[23] ;
 wire \id_ex_rs1_data[24] ;
 wire \id_ex_rs1_data[25] ;
 wire \id_ex_rs1_data[26] ;
 wire \id_ex_rs1_data[27] ;
 wire \id_ex_rs1_data[28] ;
 wire \id_ex_rs1_data[29] ;
 wire \id_ex_rs1_data[2] ;
 wire \id_ex_rs1_data[30] ;
 wire \id_ex_rs1_data[31] ;
 wire \id_ex_rs1_data[3] ;
 wire \id_ex_rs1_data[4] ;
 wire \id_ex_rs1_data[5] ;
 wire \id_ex_rs1_data[6] ;
 wire \id_ex_rs1_data[7] ;
 wire \id_ex_rs1_data[8] ;
 wire \id_ex_rs1_data[9] ;
 wire \id_ex_rs2_data[0] ;
 wire \id_ex_rs2_data[10] ;
 wire \id_ex_rs2_data[11] ;
 wire \id_ex_rs2_data[12] ;
 wire \id_ex_rs2_data[13] ;
 wire \id_ex_rs2_data[14] ;
 wire \id_ex_rs2_data[15] ;
 wire \id_ex_rs2_data[16] ;
 wire \id_ex_rs2_data[17] ;
 wire \id_ex_rs2_data[18] ;
 wire \id_ex_rs2_data[19] ;
 wire \id_ex_rs2_data[1] ;
 wire \id_ex_rs2_data[20] ;
 wire \id_ex_rs2_data[21] ;
 wire \id_ex_rs2_data[22] ;
 wire \id_ex_rs2_data[23] ;
 wire \id_ex_rs2_data[24] ;
 wire \id_ex_rs2_data[25] ;
 wire \id_ex_rs2_data[26] ;
 wire \id_ex_rs2_data[27] ;
 wire \id_ex_rs2_data[28] ;
 wire \id_ex_rs2_data[29] ;
 wire \id_ex_rs2_data[2] ;
 wire \id_ex_rs2_data[30] ;
 wire \id_ex_rs2_data[31] ;
 wire \id_ex_rs2_data[3] ;
 wire \id_ex_rs2_data[4] ;
 wire \id_ex_rs2_data[5] ;
 wire \id_ex_rs2_data[6] ;
 wire \id_ex_rs2_data[7] ;
 wire \id_ex_rs2_data[8] ;
 wire \id_ex_rs2_data[9] ;
 wire id_ex_valid;
 wire id_reg_write;
 wire if_id_valid;
 wire mem_wb_valid;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net15;
 wire net16;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \register_file.write_data[0] ;
 wire \register_file.write_data[10] ;
 wire \register_file.write_data[11] ;
 wire \register_file.write_data[12] ;
 wire \register_file.write_data[13] ;
 wire \register_file.write_data[14] ;
 wire \register_file.write_data[15] ;
 wire \register_file.write_data[16] ;
 wire \register_file.write_data[17] ;
 wire \register_file.write_data[18] ;
 wire \register_file.write_data[19] ;
 wire \register_file.write_data[1] ;
 wire \register_file.write_data[20] ;
 wire \register_file.write_data[21] ;
 wire \register_file.write_data[22] ;
 wire \register_file.write_data[23] ;
 wire \register_file.write_data[24] ;
 wire \register_file.write_data[25] ;
 wire \register_file.write_data[26] ;
 wire \register_file.write_data[27] ;
 wire \register_file.write_data[28] ;
 wire \register_file.write_data[29] ;
 wire \register_file.write_data[2] ;
 wire \register_file.write_data[30] ;
 wire \register_file.write_data[31] ;
 wire \register_file.write_data[3] ;
 wire \register_file.write_data[4] ;
 wire \register_file.write_data[5] ;
 wire \register_file.write_data[6] ;
 wire \register_file.write_data[7] ;
 wire \register_file.write_data[8] ;
 wire \register_file.write_data[9] ;

 sky130_fd_sc_hd__conb_1 CPU_core_143 (.LO(net143));
 sky130_fd_sc_hd__conb_1 CPU_core_144 (.LO(net144));
 sky130_fd_sc_hd__conb_1 CPU_core_145 (.LO(net145));
 sky130_fd_sc_hd__conb_1 CPU_core_146 (.LO(net146));
 sky130_fd_sc_hd__conb_1 CPU_core_147 (.LO(net147));
 sky130_fd_sc_hd__conb_1 CPU_core_148 (.LO(net148));
 sky130_fd_sc_hd__conb_1 CPU_core_149 (.LO(net149));
 sky130_fd_sc_hd__conb_1 CPU_core_150 (.LO(net150));
 sky130_fd_sc_hd__conb_1 CPU_core_151 (.LO(net151));
 sky130_fd_sc_hd__conb_1 CPU_core_152 (.LO(net152));
 sky130_fd_sc_hd__conb_1 CPU_core_153 (.LO(net153));
 sky130_fd_sc_hd__conb_1 CPU_core_154 (.LO(net154));
 sky130_fd_sc_hd__conb_1 CPU_core_155 (.LO(net155));
 sky130_fd_sc_hd__conb_1 CPU_core_156 (.LO(net156));
 sky130_fd_sc_hd__conb_1 CPU_core_157 (.LO(net157));
 sky130_fd_sc_hd__conb_1 CPU_core_158 (.LO(net158));
 sky130_fd_sc_hd__conb_1 CPU_core_159 (.LO(net159));
 sky130_fd_sc_hd__conb_1 CPU_core_160 (.LO(net160));
 sky130_fd_sc_hd__conb_1 CPU_core_161 (.LO(net161));
 sky130_fd_sc_hd__conb_1 CPU_core_162 (.LO(net162));
 sky130_fd_sc_hd__conb_1 CPU_core_163 (.LO(net163));
 sky130_fd_sc_hd__conb_1 CPU_core_164 (.LO(net164));
 sky130_fd_sc_hd__conb_1 CPU_core_165 (.LO(net165));
 sky130_fd_sc_hd__conb_1 CPU_core_166 (.HI(net166));
 sky130_fd_sc_hd__conb_1 CPU_core_167 (.HI(net167));
 sky130_fd_sc_hd__conb_1 CPU_core_168 (.HI(net168));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Left_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Left_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Left_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Left_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Left_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Left_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Left_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_421 ();
 sky130_fd_sc_hd__inv_2 _0842_ (.A(reset),
    .Y(_0519_));
 sky130_fd_sc_hd__buf_1 _0843_ (.A(_0519_),
    .X(_0000_));
 sky130_fd_sc_hd__buf_1 _0844_ (.A(_0519_),
    .X(_0520_));
 sky130_fd_sc_hd__and2_1 _0845_ (.A(net424),
    .B(_0520_),
    .X(_0001_));
 sky130_fd_sc_hd__buf_1 _0846_ (.A(reset),
    .X(_0521_));
 sky130_fd_sc_hd__buf_1 _0847_ (.A(_0521_),
    .X(_0522_));
 sky130_fd_sc_hd__inv_2 _0848_ (.A(net411),
    .Y(_0523_));
 sky130_fd_sc_hd__nor2_1 _0849_ (.A(_0522_),
    .B(_0523_),
    .Y(_0002_));
 sky130_fd_sc_hd__and2_1 _0850_ (.A(_0000_),
    .B(net422),
    .X(_0003_));
 sky130_fd_sc_hd__and2_1 _0851_ (.A(_0000_),
    .B(net436),
    .X(_0004_));
 sky130_fd_sc_hd__and2_1 _0852_ (.A(_0000_),
    .B(net230),
    .X(_0005_));
 sky130_fd_sc_hd__and2_1 _0853_ (.A(_0000_),
    .B(net432),
    .X(_0006_));
 sky130_fd_sc_hd__and2_1 _0854_ (.A(_0000_),
    .B(net196),
    .X(_0007_));
 sky130_fd_sc_hd__and2_1 _0855_ (.A(_0000_),
    .B(net198),
    .X(_0008_));
 sky130_fd_sc_hd__and2_1 _0856_ (.A(_0000_),
    .B(net423),
    .X(_0009_));
 sky130_fd_sc_hd__and2_1 _0857_ (.A(_0000_),
    .B(net425),
    .X(_0010_));
 sky130_fd_sc_hd__and2_1 _0858_ (.A(_0000_),
    .B(net420),
    .X(_0011_));
 sky130_fd_sc_hd__and2_1 _0859_ (.A(_0000_),
    .B(net414),
    .X(_0012_));
 sky130_fd_sc_hd__and2_1 _0860_ (.A(_0000_),
    .B(net438),
    .X(_0013_));
 sky130_fd_sc_hd__buf_1 _0861_ (.A(_0519_),
    .X(_0524_));
 sky130_fd_sc_hd__and2_1 _0862_ (.A(_0524_),
    .B(net439),
    .X(_0014_));
 sky130_fd_sc_hd__and2_1 _0863_ (.A(_0524_),
    .B(net382),
    .X(_0015_));
 sky130_fd_sc_hd__and2_1 _0864_ (.A(_0524_),
    .B(net385),
    .X(_0016_));
 sky130_fd_sc_hd__and2_1 _0865_ (.A(_0524_),
    .B(net376),
    .X(_0017_));
 sky130_fd_sc_hd__and2_1 _0866_ (.A(_0524_),
    .B(net374),
    .X(_0018_));
 sky130_fd_sc_hd__and2_1 _0867_ (.A(_0524_),
    .B(net380),
    .X(_0019_));
 sky130_fd_sc_hd__and2_1 _0868_ (.A(_0524_),
    .B(net370),
    .X(_0020_));
 sky130_fd_sc_hd__and2_1 _0869_ (.A(_0524_),
    .B(net335),
    .X(_0021_));
 sky130_fd_sc_hd__and2_1 _0870_ (.A(_0524_),
    .B(net322),
    .X(_0022_));
 sky130_fd_sc_hd__and2_1 _0871_ (.A(_0524_),
    .B(net326),
    .X(_0023_));
 sky130_fd_sc_hd__and2_1 _0872_ (.A(_0524_),
    .B(net328),
    .X(_0024_));
 sky130_fd_sc_hd__and2_1 _0873_ (.A(_0524_),
    .B(net430),
    .X(_0025_));
 sky130_fd_sc_hd__buf_1 _0874_ (.A(_0519_),
    .X(_0525_));
 sky130_fd_sc_hd__and2_1 _0875_ (.A(_0525_),
    .B(net421),
    .X(_0026_));
 sky130_fd_sc_hd__and2_1 _0876_ (.A(_0525_),
    .B(net324),
    .X(_0027_));
 sky130_fd_sc_hd__and2_1 _0877_ (.A(_0525_),
    .B(net200),
    .X(_0028_));
 sky130_fd_sc_hd__and2_1 _0878_ (.A(_0525_),
    .B(net435),
    .X(_0029_));
 sky130_fd_sc_hd__and2_1 _0879_ (.A(_0525_),
    .B(net437),
    .X(_0030_));
 sky130_fd_sc_hd__and2_1 _0880_ (.A(_0525_),
    .B(net418),
    .X(_0031_));
 sky130_fd_sc_hd__and2_1 _0881_ (.A(_0525_),
    .B(net429),
    .X(_0032_));
 sky130_fd_sc_hd__o21ai_4 _0882_ (.A1(net313),
    .A2(net308),
    .B1(net386),
    .Y(_0526_));
 sky130_fd_sc_hd__or3b_1 _0883_ (.A(net308),
    .B(_0526_),
    .C_N(\forwarding_unit.rs1_ex[0] ),
    .X(_0527_));
 sky130_fd_sc_hd__clkbuf_4 _0884_ (.A(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__mux2_1 _0885_ (.A0(\register_file.write_data[0] ),
    .A1(\id_ex_rs1_data[0] ),
    .S(_0528_),
    .X(_0529_));
 sky130_fd_sc_hd__o21ai_1 _0886_ (.A1(\forwarding_unit.rd_mem[0] ),
    .A2(\forwarding_unit.rd_mem[1] ),
    .B1(\forwarding_unit.reg_write_mem ),
    .Y(_0530_));
 sky130_fd_sc_hd__or3b_1 _0887_ (.A(_0530_),
    .B(net459),
    .C_N(\forwarding_unit.rs1_ex[0] ),
    .X(_0531_));
 sky130_fd_sc_hd__clkbuf_4 _0888_ (.A(_0531_),
    .X(_0532_));
 sky130_fd_sc_hd__mux2_1 _0889_ (.A0(net424),
    .A1(_0529_),
    .S(_0532_),
    .X(_0533_));
 sky130_fd_sc_hd__and2_1 _0890_ (.A(net506),
    .B(net395),
    .X(_0534_));
 sky130_fd_sc_hd__o21a_1 _0891_ (.A1(\forwarding_unit.rd_mem[0] ),
    .A2(\forwarding_unit.rd_mem[1] ),
    .B1(net433),
    .X(_0535_));
 sky130_fd_sc_hd__nor4b_1 _0892_ (.A(\forwarding_unit.rd_mem[0] ),
    .B(\forwarding_unit.rs2_ex[3] ),
    .C(\forwarding_unit.rs2_ex[0] ),
    .D_N(\forwarding_unit.rs2_ex[1] ),
    .Y(_0536_));
 sky130_fd_sc_hd__nand2_2 _0893_ (.A(_0535_),
    .B(net142),
    .Y(_0537_));
 sky130_fd_sc_hd__o21a_2 _0894_ (.A1(net313),
    .A2(net308),
    .B1(net386),
    .X(_0538_));
 sky130_fd_sc_hd__nor4b_1 _0895_ (.A(net313),
    .B(\forwarding_unit.rs2_ex[3] ),
    .C(\forwarding_unit.rs2_ex[0] ),
    .D_N(\forwarding_unit.rs2_ex[1] ),
    .Y(_0539_));
 sky130_fd_sc_hd__a32o_1 _0896_ (.A1(\register_file.write_data[0] ),
    .A2(_0538_),
    .A3(net141),
    .B1(_0535_),
    .B2(net543),
    .X(_0540_));
 sky130_fd_sc_hd__or4b_2 _0897_ (.A(\forwarding_unit.rd_wb[0] ),
    .B(\forwarding_unit.rs2_ex[3] ),
    .C(\forwarding_unit.rs2_ex[0] ),
    .D_N(\forwarding_unit.rs2_ex[1] ),
    .X(_0541_));
 sky130_fd_sc_hd__o21a_1 _0898_ (.A1(_0526_),
    .A2(_0541_),
    .B1(\id_ex_rs2_data[0] ),
    .X(_0542_));
 sky130_fd_sc_hd__inv_2 _0899_ (.A(net395),
    .Y(_0543_));
 sky130_fd_sc_hd__o221a_1 _0900_ (.A1(net424),
    .A2(_0537_),
    .B1(_0540_),
    .B2(_0542_),
    .C1(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__or2_1 _0901_ (.A(_0534_),
    .B(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__or2b_1 _0902_ (.A(_0533_),
    .B_N(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__or2b_1 _0903_ (.A(net507),
    .B_N(_0533_),
    .X(_0547_));
 sky130_fd_sc_hd__a21oi_1 _0904_ (.A1(_0546_),
    .A2(net508),
    .B1(_0522_),
    .Y(_0033_));
 sky130_fd_sc_hd__or2_1 _0905_ (.A(_0543_),
    .B(net526),
    .X(_0548_));
 sky130_fd_sc_hd__or3_1 _0906_ (.A(\register_file.write_data[1] ),
    .B(_0526_),
    .C(_0541_),
    .X(_0549_));
 sky130_fd_sc_hd__a21o_1 _0907_ (.A1(_0538_),
    .A2(net141),
    .B1(\id_ex_rs2_data[1] ),
    .X(_0550_));
 sky130_fd_sc_hd__a31o_1 _0908_ (.A1(\ex_mem_alu_result[1] ),
    .A2(_0535_),
    .A3(net142),
    .B1(net395),
    .X(_0551_));
 sky130_fd_sc_hd__a31o_1 _0909_ (.A1(_0537_),
    .A2(_0549_),
    .A3(_0550_),
    .B1(_0551_),
    .X(_0552_));
 sky130_fd_sc_hd__a211o_1 _0910_ (.A1(_0548_),
    .A2(_0552_),
    .B1(_0534_),
    .C1(_0544_),
    .X(_0553_));
 sky130_fd_sc_hd__o211ai_1 _0911_ (.A1(_0534_),
    .A2(_0544_),
    .B1(_0548_),
    .C1(_0552_),
    .Y(_0554_));
 sky130_fd_sc_hd__and3b_1 _0912_ (.A_N(\forwarding_unit.rd_mem[1] ),
    .B(\forwarding_unit.rs1_ex[0] ),
    .C(_0535_),
    .X(_0555_));
 sky130_fd_sc_hd__buf_2 _0913_ (.A(_0555_),
    .X(_0556_));
 sky130_fd_sc_hd__nand2_1 _0914_ (.A(net530),
    .B(_0528_),
    .Y(_0557_));
 sky130_fd_sc_hd__and3b_2 _0915_ (.A_N(\forwarding_unit.rd_wb[1] ),
    .B(_0538_),
    .C(\forwarding_unit.rs1_ex[0] ),
    .X(_0558_));
 sky130_fd_sc_hd__a21oi_1 _0916_ (.A1(\register_file.write_data[1] ),
    .A2(_0558_),
    .B1(_0556_),
    .Y(_0559_));
 sky130_fd_sc_hd__a22o_1 _0917_ (.A1(_0523_),
    .A2(_0556_),
    .B1(_0557_),
    .B2(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__a21oi_1 _0918_ (.A1(_0553_),
    .A2(_0554_),
    .B1(net531),
    .Y(_0561_));
 sky130_fd_sc_hd__nand3_1 _0919_ (.A(_0553_),
    .B(_0554_),
    .C(_0560_),
    .Y(_0562_));
 sky130_fd_sc_hd__and2b_1 _0920_ (.A_N(_0561_),
    .B(net527),
    .X(_0563_));
 sky130_fd_sc_hd__buf_1 _0921_ (.A(_0521_),
    .X(_0564_));
 sky130_fd_sc_hd__a21oi_1 _0922_ (.A1(_0546_),
    .A2(_0563_),
    .B1(_0564_),
    .Y(_0565_));
 sky130_fd_sc_hd__o21a_1 _0923_ (.A1(_0546_),
    .A2(net528),
    .B1(_0565_),
    .X(_0034_));
 sky130_fd_sc_hd__nand2_2 _0924_ (.A(_0538_),
    .B(net141),
    .Y(_0566_));
 sky130_fd_sc_hd__or4b_1 _0925_ (.A(\forwarding_unit.rd_mem[0] ),
    .B(\forwarding_unit.rs2_ex[3] ),
    .C(\forwarding_unit.rs2_ex[0] ),
    .D_N(\forwarding_unit.rs2_ex[1] ),
    .X(_0567_));
 sky130_fd_sc_hd__nor2_1 _0926_ (.A(_0530_),
    .B(_0567_),
    .Y(_0568_));
 sky130_fd_sc_hd__and3_1 _0927_ (.A(\register_file.write_data[2] ),
    .B(_0538_),
    .C(net141),
    .X(_0569_));
 sky130_fd_sc_hd__a211o_1 _0928_ (.A1(\id_ex_rs2_data[2] ),
    .A2(_0566_),
    .B1(_0568_),
    .C1(_0569_),
    .X(_0570_));
 sky130_fd_sc_hd__or2_1 _0929_ (.A(\dmem.address[2] ),
    .B(_0537_),
    .X(_0571_));
 sky130_fd_sc_hd__a31o_1 _0930_ (.A1(_0543_),
    .A2(_0570_),
    .A3(_0571_),
    .B1(_0534_),
    .X(_0572_));
 sky130_fd_sc_hd__xor2_1 _0931_ (.A(_0553_),
    .B(_0572_),
    .X(_0573_));
 sky130_fd_sc_hd__mux2_1 _0932_ (.A0(\register_file.write_data[2] ),
    .A1(\id_ex_rs1_data[2] ),
    .S(_0528_),
    .X(_0574_));
 sky130_fd_sc_hd__mux2_1 _0933_ (.A0(net422),
    .A1(_0574_),
    .S(_0532_),
    .X(_0575_));
 sky130_fd_sc_hd__xnor2_1 _0934_ (.A(_0573_),
    .B(_0575_),
    .Y(_0576_));
 sky130_fd_sc_hd__a21o_1 _0935_ (.A1(_0546_),
    .A2(net527),
    .B1(_0561_),
    .X(_0577_));
 sky130_fd_sc_hd__a21oi_1 _0936_ (.A1(_0576_),
    .A2(_0577_),
    .B1(_0564_),
    .Y(_0578_));
 sky130_fd_sc_hd__o21a_1 _0937_ (.A1(_0576_),
    .A2(_0577_),
    .B1(_0578_),
    .X(_0035_));
 sky130_fd_sc_hd__a21o_1 _0938_ (.A1(_0538_),
    .A2(net141),
    .B1(\id_ex_rs2_data[3] ),
    .X(_0579_));
 sky130_fd_sc_hd__o211a_1 _0939_ (.A1(\register_file.write_data[3] ),
    .A2(_0566_),
    .B1(_0537_),
    .C1(_0579_),
    .X(_0580_));
 sky130_fd_sc_hd__a31o_1 _0940_ (.A1(\dmem.address[3] ),
    .A2(_0535_),
    .A3(net142),
    .B1(net395),
    .X(_0581_));
 sky130_fd_sc_hd__o22a_1 _0941_ (.A1(_0543_),
    .A2(net520),
    .B1(_0580_),
    .B2(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__or3_1 _0942_ (.A(_0553_),
    .B(_0572_),
    .C(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__buf_2 _0943_ (.A(_0583_),
    .X(_0584_));
 sky130_fd_sc_hd__o21ai_1 _0944_ (.A1(_0553_),
    .A2(_0572_),
    .B1(_0582_),
    .Y(_0585_));
 sky130_fd_sc_hd__nand2_1 _0945_ (.A(_0584_),
    .B(net521),
    .Y(_0586_));
 sky130_fd_sc_hd__mux2_1 _0946_ (.A0(\register_file.write_data[3] ),
    .A1(\id_ex_rs1_data[3] ),
    .S(_0528_),
    .X(_0587_));
 sky130_fd_sc_hd__mux2_1 _0947_ (.A0(net436),
    .A1(_0587_),
    .S(_0532_),
    .X(_0588_));
 sky130_fd_sc_hd__xnor2_1 _0948_ (.A(_0586_),
    .B(_0588_),
    .Y(_0589_));
 sky130_fd_sc_hd__and2b_1 _0949_ (.A_N(_0573_),
    .B(_0575_),
    .X(_0590_));
 sky130_fd_sc_hd__a21oi_1 _0950_ (.A1(_0576_),
    .A2(_0577_),
    .B1(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__buf_1 _0951_ (.A(_0519_),
    .X(_0592_));
 sky130_fd_sc_hd__o21ai_1 _0952_ (.A1(net522),
    .A2(_0591_),
    .B1(_0592_),
    .Y(_0593_));
 sky130_fd_sc_hd__a21oi_1 _0953_ (.A1(net522),
    .A2(_0591_),
    .B1(_0593_),
    .Y(_0036_));
 sky130_fd_sc_hd__clkbuf_4 _0954_ (.A(_0568_),
    .X(_0594_));
 sky130_fd_sc_hd__mux2_1 _0955_ (.A0(\register_file.write_data[4] ),
    .A1(\id_ex_rs2_data[4] ),
    .S(_0566_),
    .X(_0595_));
 sky130_fd_sc_hd__or2_1 _0956_ (.A(net230),
    .B(_0537_),
    .X(_0596_));
 sky130_fd_sc_hd__o211a_1 _0957_ (.A1(_0594_),
    .A2(_0595_),
    .B1(_0596_),
    .C1(_0543_),
    .X(_0597_));
 sky130_fd_sc_hd__xnor2_1 _0958_ (.A(_0584_),
    .B(net396),
    .Y(_0598_));
 sky130_fd_sc_hd__mux2_1 _0959_ (.A0(\register_file.write_data[4] ),
    .A1(\id_ex_rs1_data[4] ),
    .S(_0528_),
    .X(_0599_));
 sky130_fd_sc_hd__mux2_1 _0960_ (.A0(net230),
    .A1(_0599_),
    .S(_0532_),
    .X(_0600_));
 sky130_fd_sc_hd__nand2_1 _0961_ (.A(net397),
    .B(_0600_),
    .Y(_0601_));
 sky130_fd_sc_hd__or2_1 _0962_ (.A(net397),
    .B(_0600_),
    .X(_0602_));
 sky130_fd_sc_hd__nand2_1 _0963_ (.A(net398),
    .B(_0602_),
    .Y(_0603_));
 sky130_fd_sc_hd__nand2_1 _0964_ (.A(_0586_),
    .B(_0588_),
    .Y(_0604_));
 sky130_fd_sc_hd__o21a_1 _0965_ (.A1(_0589_),
    .A2(_0591_),
    .B1(_0604_),
    .X(_0605_));
 sky130_fd_sc_hd__or2_1 _0966_ (.A(_0603_),
    .B(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__buf_1 _0967_ (.A(_0521_),
    .X(_0607_));
 sky130_fd_sc_hd__a21oi_1 _0968_ (.A1(_0603_),
    .A2(_0605_),
    .B1(_0607_),
    .Y(_0608_));
 sky130_fd_sc_hd__and2_1 _0969_ (.A(_0606_),
    .B(_0608_),
    .X(_0037_));
 sky130_fd_sc_hd__buf_4 _0970_ (.A(_0566_),
    .X(_0609_));
 sky130_fd_sc_hd__mux2_1 _0971_ (.A0(\register_file.write_data[5] ),
    .A1(\id_ex_rs2_data[5] ),
    .S(_0609_),
    .X(_0610_));
 sky130_fd_sc_hd__buf_2 _0972_ (.A(_0537_),
    .X(_0611_));
 sky130_fd_sc_hd__or2_1 _0973_ (.A(\dmem.address[5] ),
    .B(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__clkbuf_4 _0974_ (.A(_0543_),
    .X(_0613_));
 sky130_fd_sc_hd__o211a_1 _0975_ (.A1(_0594_),
    .A2(_0610_),
    .B1(_0612_),
    .C1(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__or2_2 _0976_ (.A(net396),
    .B(_0614_),
    .X(_0615_));
 sky130_fd_sc_hd__nor2_1 _0977_ (.A(_0584_),
    .B(_0615_),
    .Y(_0616_));
 sky130_fd_sc_hd__o21a_1 _0978_ (.A1(_0584_),
    .A2(net396),
    .B1(_0614_),
    .X(_0617_));
 sky130_fd_sc_hd__clkbuf_4 _0979_ (.A(_0528_),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_1 _0980_ (.A0(\register_file.write_data[5] ),
    .A1(\id_ex_rs1_data[5] ),
    .S(_0618_),
    .X(_0619_));
 sky130_fd_sc_hd__buf_4 _0981_ (.A(_0532_),
    .X(_0620_));
 sky130_fd_sc_hd__mux2_1 _0982_ (.A0(\dmem.address[5] ),
    .A1(_0619_),
    .S(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__o21ai_1 _0983_ (.A1(_0616_),
    .A2(_0617_),
    .B1(_0621_),
    .Y(_0622_));
 sky130_fd_sc_hd__nor3_1 _0984_ (.A(_0616_),
    .B(_0617_),
    .C(_0621_),
    .Y(_0623_));
 sky130_fd_sc_hd__inv_2 _0985_ (.A(_0623_),
    .Y(_0624_));
 sky130_fd_sc_hd__nand2_1 _0986_ (.A(_0622_),
    .B(_0624_),
    .Y(_0625_));
 sky130_fd_sc_hd__a21oi_1 _0987_ (.A1(net398),
    .A2(_0606_),
    .B1(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hd__a31o_1 _0988_ (.A1(net398),
    .A2(_0606_),
    .A3(_0625_),
    .B1(_0607_),
    .X(_0627_));
 sky130_fd_sc_hd__nor2_1 _0989_ (.A(net399),
    .B(_0627_),
    .Y(_0038_));
 sky130_fd_sc_hd__buf_1 _0990_ (.A(_0519_),
    .X(_0628_));
 sky130_fd_sc_hd__mux2_1 _0991_ (.A0(\register_file.write_data[6] ),
    .A1(\id_ex_rs2_data[6] ),
    .S(_0566_),
    .X(_0629_));
 sky130_fd_sc_hd__or2_1 _0992_ (.A(\dmem.address[6] ),
    .B(_0537_),
    .X(_0630_));
 sky130_fd_sc_hd__o211a_1 _0993_ (.A1(_0594_),
    .A2(_0629_),
    .B1(_0630_),
    .C1(_0543_),
    .X(_0631_));
 sky130_fd_sc_hd__xnor2_1 _0994_ (.A(_0616_),
    .B(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hd__mux2_1 _0995_ (.A0(\register_file.write_data[6] ),
    .A1(\id_ex_rs1_data[6] ),
    .S(_0618_),
    .X(_0633_));
 sky130_fd_sc_hd__mux2_1 _0996_ (.A0(net196),
    .A1(_0633_),
    .S(_0620_),
    .X(_0634_));
 sky130_fd_sc_hd__or2b_1 _0997_ (.A(_0632_),
    .B_N(_0634_),
    .X(_0635_));
 sky130_fd_sc_hd__or2b_1 _0998_ (.A(_0634_),
    .B_N(_0632_),
    .X(_0636_));
 sky130_fd_sc_hd__nand2_1 _0999_ (.A(_0635_),
    .B(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__o211a_1 _1000_ (.A1(_0603_),
    .A2(_0605_),
    .B1(_0622_),
    .C1(_0601_),
    .X(_0638_));
 sky130_fd_sc_hd__or2_1 _1001_ (.A(net139),
    .B(_0638_),
    .X(_0639_));
 sky130_fd_sc_hd__nand2_1 _1002_ (.A(_0637_),
    .B(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__or2_1 _1003_ (.A(_0637_),
    .B(_0639_),
    .X(_0641_));
 sky130_fd_sc_hd__and3_1 _1004_ (.A(_0628_),
    .B(_0640_),
    .C(_0641_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _1005_ (.A0(\register_file.write_data[7] ),
    .A1(\id_ex_rs2_data[7] ),
    .S(_0566_),
    .X(_0642_));
 sky130_fd_sc_hd__or2_1 _1006_ (.A(\dmem.address[7] ),
    .B(_0537_),
    .X(_0643_));
 sky130_fd_sc_hd__o211a_1 _1007_ (.A1(_0594_),
    .A2(_0642_),
    .B1(_0643_),
    .C1(_0543_),
    .X(_0644_));
 sky130_fd_sc_hd__or2_1 _1008_ (.A(_0631_),
    .B(_0644_),
    .X(_0645_));
 sky130_fd_sc_hd__nor3_2 _1009_ (.A(_0584_),
    .B(_0615_),
    .C(_0645_),
    .Y(_0646_));
 sky130_fd_sc_hd__o31a_1 _1010_ (.A1(_0584_),
    .A2(_0615_),
    .A3(_0631_),
    .B1(_0644_),
    .X(_0647_));
 sky130_fd_sc_hd__or2_1 _1011_ (.A(_0646_),
    .B(_0647_),
    .X(_0648_));
 sky130_fd_sc_hd__mux2_1 _1012_ (.A0(\register_file.write_data[7] ),
    .A1(\id_ex_rs1_data[7] ),
    .S(_0528_),
    .X(_0649_));
 sky130_fd_sc_hd__mux2_1 _1013_ (.A0(net198),
    .A1(_0649_),
    .S(_0532_),
    .X(_0650_));
 sky130_fd_sc_hd__nand2_1 _1014_ (.A(_0648_),
    .B(_0650_),
    .Y(_0651_));
 sky130_fd_sc_hd__or3_1 _1015_ (.A(_0646_),
    .B(_0647_),
    .C(_0650_),
    .X(_0652_));
 sky130_fd_sc_hd__nand2_1 _1016_ (.A(_0651_),
    .B(_0652_),
    .Y(_0653_));
 sky130_fd_sc_hd__a21oi_1 _1017_ (.A1(_0635_),
    .A2(_0641_),
    .B1(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__a31o_1 _1018_ (.A1(_0635_),
    .A2(_0641_),
    .A3(_0653_),
    .B1(_0607_),
    .X(_0655_));
 sky130_fd_sc_hd__nor2_1 _1019_ (.A(_0654_),
    .B(_0655_),
    .Y(_0040_));
 sky130_fd_sc_hd__and3b_1 _1020_ (.A_N(_0632_),
    .B(_0634_),
    .C(_0652_),
    .X(_0656_));
 sky130_fd_sc_hd__a21oi_1 _1021_ (.A1(_0648_),
    .A2(_0650_),
    .B1(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__o41a_2 _1022_ (.A1(net139),
    .A2(_0637_),
    .A3(_0638_),
    .A4(_0653_),
    .B1(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__or3_1 _1023_ (.A(_0584_),
    .B(_0615_),
    .C(_0645_),
    .X(_0659_));
 sky130_fd_sc_hd__buf_2 _1024_ (.A(_0659_),
    .X(_0660_));
 sky130_fd_sc_hd__and3_1 _1025_ (.A(\register_file.write_data[8] ),
    .B(_0538_),
    .C(net542),
    .X(_0661_));
 sky130_fd_sc_hd__o21a_1 _1026_ (.A1(_0526_),
    .A2(_0541_),
    .B1(\id_ex_rs2_data[8] ),
    .X(_0662_));
 sky130_fd_sc_hd__or3_1 _1027_ (.A(\dmem.address[8] ),
    .B(_0530_),
    .C(_0567_),
    .X(_0663_));
 sky130_fd_sc_hd__o311a_1 _1028_ (.A1(_0568_),
    .A2(_0661_),
    .A3(_0662_),
    .B1(_0663_),
    .C1(_0543_),
    .X(_0664_));
 sky130_fd_sc_hd__xnor2_1 _1029_ (.A(_0660_),
    .B(_0664_),
    .Y(_0665_));
 sky130_fd_sc_hd__mux2_1 _1030_ (.A0(\register_file.write_data[8] ),
    .A1(\id_ex_rs1_data[8] ),
    .S(_0618_),
    .X(_0666_));
 sky130_fd_sc_hd__mux2_1 _1031_ (.A0(net423),
    .A1(_0666_),
    .S(_0620_),
    .X(_0667_));
 sky130_fd_sc_hd__xnor2_1 _1032_ (.A(_0665_),
    .B(_0667_),
    .Y(_0668_));
 sky130_fd_sc_hd__nand2_1 _1033_ (.A(_0658_),
    .B(_0668_),
    .Y(_0669_));
 sky130_fd_sc_hd__or2_1 _1034_ (.A(_0658_),
    .B(_0668_),
    .X(_0670_));
 sky130_fd_sc_hd__and3_1 _1035_ (.A(_0628_),
    .B(_0669_),
    .C(_0670_),
    .X(_0041_));
 sky130_fd_sc_hd__nand2_1 _1036_ (.A(_0665_),
    .B(_0667_),
    .Y(_0671_));
 sky130_fd_sc_hd__or4_1 _1037_ (.A(_0584_),
    .B(_0615_),
    .C(_0645_),
    .D(_0664_),
    .X(_0672_));
 sky130_fd_sc_hd__and3_1 _1038_ (.A(\register_file.write_data[9] ),
    .B(_0538_),
    .C(net542),
    .X(_0673_));
 sky130_fd_sc_hd__o21a_1 _1039_ (.A1(_0526_),
    .A2(_0541_),
    .B1(\id_ex_rs2_data[9] ),
    .X(_0674_));
 sky130_fd_sc_hd__or3_1 _1040_ (.A(\dmem.address[9] ),
    .B(_0530_),
    .C(_0567_),
    .X(_0675_));
 sky130_fd_sc_hd__o311a_1 _1041_ (.A1(_0568_),
    .A2(_0673_),
    .A3(_0674_),
    .B1(_0675_),
    .C1(_0543_),
    .X(_0676_));
 sky130_fd_sc_hd__xnor2_1 _1042_ (.A(_0672_),
    .B(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__mux2_1 _1043_ (.A0(\register_file.write_data[9] ),
    .A1(\id_ex_rs1_data[9] ),
    .S(_0618_),
    .X(_0678_));
 sky130_fd_sc_hd__mux2_1 _1044_ (.A0(net425),
    .A1(_0678_),
    .S(_0620_),
    .X(_0679_));
 sky130_fd_sc_hd__xnor2_1 _1045_ (.A(_0677_),
    .B(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__a21oi_1 _1046_ (.A1(_0671_),
    .A2(_0670_),
    .B1(_0680_),
    .Y(_0681_));
 sky130_fd_sc_hd__a31o_1 _1047_ (.A1(_0671_),
    .A2(_0670_),
    .A3(_0680_),
    .B1(_0607_),
    .X(_0682_));
 sky130_fd_sc_hd__nor2_1 _1048_ (.A(_0681_),
    .B(_0682_),
    .Y(_0042_));
 sky130_fd_sc_hd__or2_1 _1049_ (.A(_0664_),
    .B(_0676_),
    .X(_0683_));
 sky130_fd_sc_hd__mux2_1 _1050_ (.A0(\register_file.write_data[10] ),
    .A1(\id_ex_rs2_data[10] ),
    .S(_0609_),
    .X(_0684_));
 sky130_fd_sc_hd__or2_1 _1051_ (.A(\dmem.address[10] ),
    .B(_0611_),
    .X(_0685_));
 sky130_fd_sc_hd__o211a_1 _1052_ (.A1(_0594_),
    .A2(_0684_),
    .B1(_0685_),
    .C1(_0613_),
    .X(_0686_));
 sky130_fd_sc_hd__or2_1 _1053_ (.A(_0683_),
    .B(_0686_),
    .X(_0687_));
 sky130_fd_sc_hd__o21ai_1 _1054_ (.A1(_0660_),
    .A2(_0683_),
    .B1(_0686_),
    .Y(_0688_));
 sky130_fd_sc_hd__o21ai_2 _1055_ (.A1(_0660_),
    .A2(_0687_),
    .B1(_0688_),
    .Y(_0689_));
 sky130_fd_sc_hd__buf_4 _1056_ (.A(_0618_),
    .X(_0690_));
 sky130_fd_sc_hd__mux2_1 _1057_ (.A0(net538),
    .A1(\id_ex_rs1_data[10] ),
    .S(_0690_),
    .X(_0691_));
 sky130_fd_sc_hd__buf_4 _1058_ (.A(_0620_),
    .X(_0692_));
 sky130_fd_sc_hd__mux2_1 _1059_ (.A0(net420),
    .A1(_0691_),
    .S(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__xor2_2 _1060_ (.A(_0689_),
    .B(_0693_),
    .X(_0694_));
 sky130_fd_sc_hd__nor2_1 _1061_ (.A(_0677_),
    .B(_0679_),
    .Y(_0695_));
 sky130_fd_sc_hd__nand2_1 _1062_ (.A(_0677_),
    .B(_0679_),
    .Y(_0696_));
 sky130_fd_sc_hd__o21ai_1 _1063_ (.A1(_0671_),
    .A2(_0695_),
    .B1(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__nor2_1 _1064_ (.A(_0668_),
    .B(_0680_),
    .Y(_0698_));
 sky130_fd_sc_hd__and2b_1 _1065_ (.A_N(_0658_),
    .B(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__or2_1 _1066_ (.A(_0697_),
    .B(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__or2_1 _1067_ (.A(_0694_),
    .B(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__nand2_1 _1068_ (.A(_0694_),
    .B(_0700_),
    .Y(_0702_));
 sky130_fd_sc_hd__and3_1 _1069_ (.A(_0628_),
    .B(_0701_),
    .C(_0702_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _1070_ (.A0(\register_file.write_data[11] ),
    .A1(\id_ex_rs2_data[11] ),
    .S(_0609_),
    .X(_0703_));
 sky130_fd_sc_hd__or2_1 _1071_ (.A(\dmem.address[11] ),
    .B(_0611_),
    .X(_0704_));
 sky130_fd_sc_hd__o211a_1 _1072_ (.A1(_0594_),
    .A2(_0703_),
    .B1(_0704_),
    .C1(_0613_),
    .X(_0705_));
 sky130_fd_sc_hd__or2_1 _1073_ (.A(_0687_),
    .B(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__nor2_1 _1074_ (.A(_0660_),
    .B(_0706_),
    .Y(_0707_));
 sky130_fd_sc_hd__o21a_1 _1075_ (.A1(_0660_),
    .A2(_0687_),
    .B1(_0705_),
    .X(_0708_));
 sky130_fd_sc_hd__mux2_1 _1076_ (.A0(\register_file.write_data[11] ),
    .A1(\id_ex_rs1_data[11] ),
    .S(_0528_),
    .X(_0709_));
 sky130_fd_sc_hd__mux2_1 _1077_ (.A0(net414),
    .A1(_0709_),
    .S(_0532_),
    .X(_0710_));
 sky130_fd_sc_hd__o21ai_1 _1078_ (.A1(_0707_),
    .A2(_0708_),
    .B1(_0710_),
    .Y(_0711_));
 sky130_fd_sc_hd__or3_1 _1079_ (.A(_0707_),
    .B(_0708_),
    .C(_0710_),
    .X(_0712_));
 sky130_fd_sc_hd__and2_1 _1080_ (.A(_0711_),
    .B(_0712_),
    .X(_0713_));
 sky130_fd_sc_hd__a21bo_1 _1081_ (.A1(_0689_),
    .A2(_0693_),
    .B1_N(_0702_),
    .X(_0714_));
 sky130_fd_sc_hd__a21o_1 _1082_ (.A1(_0713_),
    .A2(_0714_),
    .B1(_0521_),
    .X(_0715_));
 sky130_fd_sc_hd__o21ba_1 _1083_ (.A1(_0713_),
    .A2(_0714_),
    .B1_N(_0715_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _1084_ (.A0(\register_file.write_data[12] ),
    .A1(\id_ex_rs2_data[12] ),
    .S(_0609_),
    .X(_0716_));
 sky130_fd_sc_hd__o21a_1 _1085_ (.A1(\dmem.address[12] ),
    .A2(_0611_),
    .B1(_0613_),
    .X(_0717_));
 sky130_fd_sc_hd__o21ai_2 _1086_ (.A1(_0594_),
    .A2(_0716_),
    .B1(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hd__or3b_1 _1087_ (.A(_0660_),
    .B(_0706_),
    .C_N(_0718_),
    .X(_0719_));
 sky130_fd_sc_hd__nor2_1 _1088_ (.A(_0687_),
    .B(_0705_),
    .Y(_0720_));
 sky130_fd_sc_hd__a21o_1 _1089_ (.A1(_0646_),
    .A2(_0720_),
    .B1(_0718_),
    .X(_0721_));
 sky130_fd_sc_hd__or2_1 _1090_ (.A(\register_file.write_data[12] ),
    .B(_0618_),
    .X(_0722_));
 sky130_fd_sc_hd__o211a_1 _1091_ (.A1(\id_ex_rs1_data[12] ),
    .A2(_0558_),
    .B1(_0722_),
    .C1(_0620_),
    .X(_0723_));
 sky130_fd_sc_hd__a21oi_1 _1092_ (.A1(net438),
    .A2(_0556_),
    .B1(_0723_),
    .Y(_0724_));
 sky130_fd_sc_hd__a21o_1 _1093_ (.A1(_0719_),
    .A2(_0721_),
    .B1(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__nand3_1 _1094_ (.A(_0719_),
    .B(_0721_),
    .C(_0724_),
    .Y(_0726_));
 sky130_fd_sc_hd__nand2_1 _1095_ (.A(_0725_),
    .B(_0726_),
    .Y(_0727_));
 sky130_fd_sc_hd__nand4_1 _1096_ (.A(_0694_),
    .B(_0698_),
    .C(_0711_),
    .D(_0712_),
    .Y(_0728_));
 sky130_fd_sc_hd__and3_1 _1097_ (.A(_0689_),
    .B(_0693_),
    .C(_0712_),
    .X(_0729_));
 sky130_fd_sc_hd__inv_2 _1098_ (.A(_0711_),
    .Y(_0730_));
 sky130_fd_sc_hd__a311oi_2 _1099_ (.A1(_0694_),
    .A2(_0697_),
    .A3(_0712_),
    .B1(_0729_),
    .C1(_0730_),
    .Y(_0731_));
 sky130_fd_sc_hd__o21a_1 _1100_ (.A1(_0658_),
    .A2(_0728_),
    .B1(_0731_),
    .X(_0732_));
 sky130_fd_sc_hd__nand2_1 _1101_ (.A(_0727_),
    .B(_0732_),
    .Y(_0733_));
 sky130_fd_sc_hd__or2_1 _1102_ (.A(_0727_),
    .B(_0732_),
    .X(_0734_));
 sky130_fd_sc_hd__and3_1 _1103_ (.A(_0628_),
    .B(_0733_),
    .C(_0734_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _1104_ (.A0(\register_file.write_data[13] ),
    .A1(\id_ex_rs2_data[13] ),
    .S(_0609_),
    .X(_0735_));
 sky130_fd_sc_hd__o21a_1 _1105_ (.A1(\dmem.address[13] ),
    .A2(_0611_),
    .B1(_0613_),
    .X(_0736_));
 sky130_fd_sc_hd__o21ai_1 _1106_ (.A1(_0594_),
    .A2(_0735_),
    .B1(_0736_),
    .Y(_0737_));
 sky130_fd_sc_hd__nand2_1 _1107_ (.A(_0718_),
    .B(_0737_),
    .Y(_0738_));
 sky130_fd_sc_hd__or3_1 _1108_ (.A(_0660_),
    .B(_0706_),
    .C(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__a31o_1 _1109_ (.A1(_0646_),
    .A2(_0720_),
    .A3(_0718_),
    .B1(_0737_),
    .X(_0740_));
 sky130_fd_sc_hd__or2_1 _1110_ (.A(\register_file.write_data[13] ),
    .B(_0528_),
    .X(_0741_));
 sky130_fd_sc_hd__o211a_1 _1111_ (.A1(\id_ex_rs1_data[13] ),
    .A2(_0558_),
    .B1(_0741_),
    .C1(_0532_),
    .X(_0742_));
 sky130_fd_sc_hd__a21oi_1 _1112_ (.A1(net439),
    .A2(_0556_),
    .B1(_0742_),
    .Y(_0743_));
 sky130_fd_sc_hd__and3_1 _1113_ (.A(_0739_),
    .B(_0740_),
    .C(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__a21o_1 _1114_ (.A1(_0739_),
    .A2(_0740_),
    .B1(_0743_),
    .X(_0745_));
 sky130_fd_sc_hd__or2b_1 _1115_ (.A(_0744_),
    .B_N(_0745_),
    .X(_0746_));
 sky130_fd_sc_hd__a21oi_1 _1116_ (.A1(_0725_),
    .A2(_0734_),
    .B1(_0746_),
    .Y(_0747_));
 sky130_fd_sc_hd__a31o_1 _1117_ (.A1(_0725_),
    .A2(_0734_),
    .A3(_0746_),
    .B1(_0607_),
    .X(_0748_));
 sky130_fd_sc_hd__nor2_1 _1118_ (.A(_0747_),
    .B(_0748_),
    .Y(_0046_));
 sky130_fd_sc_hd__mux2_1 _1119_ (.A0(\register_file.write_data[14] ),
    .A1(\id_ex_rs2_data[14] ),
    .S(_0609_),
    .X(_0749_));
 sky130_fd_sc_hd__or2_1 _1120_ (.A(\dmem.address[14] ),
    .B(_0611_),
    .X(_0750_));
 sky130_fd_sc_hd__o211a_1 _1121_ (.A1(_0594_),
    .A2(_0749_),
    .B1(_0750_),
    .C1(_0613_),
    .X(_0751_));
 sky130_fd_sc_hd__or2_1 _1122_ (.A(_0738_),
    .B(_0751_),
    .X(_0752_));
 sky130_fd_sc_hd__or3_1 _1123_ (.A(_0660_),
    .B(_0706_),
    .C(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__a21boi_1 _1124_ (.A1(_0739_),
    .A2(_0751_),
    .B1_N(_0753_),
    .Y(_0754_));
 sky130_fd_sc_hd__mux2_1 _1125_ (.A0(\register_file.write_data[14] ),
    .A1(\id_ex_rs1_data[14] ),
    .S(_0618_),
    .X(_0755_));
 sky130_fd_sc_hd__mux2_1 _1126_ (.A0(net382),
    .A1(_0755_),
    .S(_0620_),
    .X(_0756_));
 sky130_fd_sc_hd__xor2_1 _1127_ (.A(_0754_),
    .B(_0756_),
    .X(_0757_));
 sky130_fd_sc_hd__o21a_1 _1128_ (.A1(_0725_),
    .A2(_0744_),
    .B1(_0745_),
    .X(_0758_));
 sky130_fd_sc_hd__o21a_1 _1129_ (.A1(_0734_),
    .A2(_0746_),
    .B1(_0758_),
    .X(_0759_));
 sky130_fd_sc_hd__nand2_1 _1130_ (.A(_0757_),
    .B(_0759_),
    .Y(_0760_));
 sky130_fd_sc_hd__or2_1 _1131_ (.A(_0757_),
    .B(_0759_),
    .X(_0761_));
 sky130_fd_sc_hd__and3_1 _1132_ (.A(_0628_),
    .B(_0760_),
    .C(_0761_),
    .X(_0047_));
 sky130_fd_sc_hd__or2b_1 _1133_ (.A(_0754_),
    .B_N(_0756_),
    .X(_0762_));
 sky130_fd_sc_hd__mux2_1 _1134_ (.A0(\register_file.write_data[15] ),
    .A1(\id_ex_rs2_data[15] ),
    .S(_0609_),
    .X(_0763_));
 sky130_fd_sc_hd__or2_1 _1135_ (.A(\dmem.address[15] ),
    .B(_0611_),
    .X(_0764_));
 sky130_fd_sc_hd__o211a_1 _1136_ (.A1(_0594_),
    .A2(_0763_),
    .B1(_0764_),
    .C1(_0613_),
    .X(_0765_));
 sky130_fd_sc_hd__xnor2_1 _1137_ (.A(_0753_),
    .B(_0765_),
    .Y(_0766_));
 sky130_fd_sc_hd__mux2_1 _1138_ (.A0(\register_file.write_data[15] ),
    .A1(\id_ex_rs1_data[15] ),
    .S(_0618_),
    .X(_0767_));
 sky130_fd_sc_hd__mux2_1 _1139_ (.A0(net385),
    .A1(_0767_),
    .S(_0620_),
    .X(_0768_));
 sky130_fd_sc_hd__xnor2_1 _1140_ (.A(_0766_),
    .B(_0768_),
    .Y(_0769_));
 sky130_fd_sc_hd__a21oi_1 _1141_ (.A1(_0762_),
    .A2(_0761_),
    .B1(_0769_),
    .Y(_0770_));
 sky130_fd_sc_hd__a31o_1 _1142_ (.A1(_0762_),
    .A2(_0761_),
    .A3(_0769_),
    .B1(_0607_),
    .X(_0771_));
 sky130_fd_sc_hd__nor2_1 _1143_ (.A(_0770_),
    .B(_0771_),
    .Y(_0048_));
 sky130_fd_sc_hd__or4_1 _1144_ (.A(_0660_),
    .B(_0706_),
    .C(_0752_),
    .D(_0765_),
    .X(_0772_));
 sky130_fd_sc_hd__buf_2 _1145_ (.A(_0772_),
    .X(_0773_));
 sky130_fd_sc_hd__mux2_1 _1146_ (.A0(\register_file.write_data[16] ),
    .A1(\id_ex_rs2_data[16] ),
    .S(_0609_),
    .X(_0774_));
 sky130_fd_sc_hd__or2_1 _1147_ (.A(\dmem.address[16] ),
    .B(_0611_),
    .X(_0775_));
 sky130_fd_sc_hd__o211a_1 _1148_ (.A1(_0594_),
    .A2(_0774_),
    .B1(_0775_),
    .C1(_0613_),
    .X(_0776_));
 sky130_fd_sc_hd__xnor2_1 _1149_ (.A(_0773_),
    .B(_0776_),
    .Y(_0777_));
 sky130_fd_sc_hd__mux2_1 _1150_ (.A0(\register_file.write_data[16] ),
    .A1(\id_ex_rs1_data[16] ),
    .S(_0618_),
    .X(_0778_));
 sky130_fd_sc_hd__mux2_1 _1151_ (.A0(net376),
    .A1(_0778_),
    .S(_0620_),
    .X(_0779_));
 sky130_fd_sc_hd__nand2_1 _1152_ (.A(_0777_),
    .B(_0779_),
    .Y(_0780_));
 sky130_fd_sc_hd__or2_1 _1153_ (.A(_0777_),
    .B(_0779_),
    .X(_0781_));
 sky130_fd_sc_hd__nand2_1 _1154_ (.A(_0780_),
    .B(_0781_),
    .Y(_0782_));
 sky130_fd_sc_hd__or4_1 _1155_ (.A(_0727_),
    .B(_0746_),
    .C(_0757_),
    .D(_0769_),
    .X(_0783_));
 sky130_fd_sc_hd__or3_1 _1156_ (.A(_0658_),
    .B(_0728_),
    .C(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__nor2_1 _1157_ (.A(_0766_),
    .B(_0768_),
    .Y(_0785_));
 sky130_fd_sc_hd__nand2_1 _1158_ (.A(_0766_),
    .B(_0768_),
    .Y(_0786_));
 sky130_fd_sc_hd__o21a_1 _1159_ (.A1(_0762_),
    .A2(_0785_),
    .B1(_0786_),
    .X(_0787_));
 sky130_fd_sc_hd__or3_1 _1160_ (.A(_0757_),
    .B(_0758_),
    .C(_0769_),
    .X(_0788_));
 sky130_fd_sc_hd__o211a_1 _1161_ (.A1(_0731_),
    .A2(_0783_),
    .B1(_0787_),
    .C1(_0788_),
    .X(_0789_));
 sky130_fd_sc_hd__and2_1 _1162_ (.A(_0784_),
    .B(_0789_),
    .X(_0790_));
 sky130_fd_sc_hd__nand2_1 _1163_ (.A(_0782_),
    .B(_0790_),
    .Y(_0791_));
 sky130_fd_sc_hd__or2_1 _1164_ (.A(_0782_),
    .B(_0790_),
    .X(_0792_));
 sky130_fd_sc_hd__and3_1 _1165_ (.A(_0628_),
    .B(_0791_),
    .C(_0792_),
    .X(_0049_));
 sky130_fd_sc_hd__and4bb_1 _1166_ (.A_N(_0765_),
    .B_N(_0752_),
    .C(_0720_),
    .D(_0646_),
    .X(_0793_));
 sky130_fd_sc_hd__clkbuf_4 _1167_ (.A(_0594_),
    .X(_0794_));
 sky130_fd_sc_hd__mux2_1 _1168_ (.A0(\register_file.write_data[17] ),
    .A1(\id_ex_rs2_data[17] ),
    .S(_0609_),
    .X(_0795_));
 sky130_fd_sc_hd__or2_1 _1169_ (.A(\dmem.address[17] ),
    .B(_0611_),
    .X(_0796_));
 sky130_fd_sc_hd__o211a_1 _1170_ (.A1(_0794_),
    .A2(_0795_),
    .B1(_0796_),
    .C1(_0613_),
    .X(_0797_));
 sky130_fd_sc_hd__nor2_1 _1171_ (.A(_0776_),
    .B(_0797_),
    .Y(_0798_));
 sky130_fd_sc_hd__nand2_1 _1172_ (.A(_0793_),
    .B(_0798_),
    .Y(_0799_));
 sky130_fd_sc_hd__o21ai_1 _1173_ (.A1(_0773_),
    .A2(_0776_),
    .B1(_0797_),
    .Y(_0800_));
 sky130_fd_sc_hd__or2_1 _1174_ (.A(\register_file.write_data[17] ),
    .B(_0618_),
    .X(_0801_));
 sky130_fd_sc_hd__o211a_1 _1175_ (.A1(\id_ex_rs1_data[17] ),
    .A2(_0558_),
    .B1(_0801_),
    .C1(_0620_),
    .X(_0802_));
 sky130_fd_sc_hd__a21oi_1 _1176_ (.A1(net374),
    .A2(_0556_),
    .B1(_0802_),
    .Y(_0803_));
 sky130_fd_sc_hd__and3_1 _1177_ (.A(_0799_),
    .B(_0800_),
    .C(_0803_),
    .X(_0804_));
 sky130_fd_sc_hd__a21o_1 _1178_ (.A1(_0799_),
    .A2(_0800_),
    .B1(_0803_),
    .X(_0805_));
 sky130_fd_sc_hd__or2b_1 _1179_ (.A(_0804_),
    .B_N(_0805_),
    .X(_0806_));
 sky130_fd_sc_hd__a21oi_1 _1180_ (.A1(_0780_),
    .A2(_0792_),
    .B1(_0806_),
    .Y(_0807_));
 sky130_fd_sc_hd__a31o_1 _1181_ (.A1(_0780_),
    .A2(_0792_),
    .A3(_0806_),
    .B1(_0607_),
    .X(_0808_));
 sky130_fd_sc_hd__nor2_1 _1182_ (.A(_0807_),
    .B(_0808_),
    .Y(_0050_));
 sky130_fd_sc_hd__mux2_1 _1183_ (.A0(\register_file.write_data[18] ),
    .A1(\id_ex_rs2_data[18] ),
    .S(_0609_),
    .X(_0809_));
 sky130_fd_sc_hd__mux2_1 _1184_ (.A0(\dmem.address[18] ),
    .A1(_0809_),
    .S(_0611_),
    .X(_0810_));
 sky130_fd_sc_hd__nand2_1 _1185_ (.A(_0613_),
    .B(_0810_),
    .Y(_0811_));
 sky130_fd_sc_hd__nand2_1 _1186_ (.A(_0798_),
    .B(_0811_),
    .Y(_0812_));
 sky130_fd_sc_hd__nor2_1 _1187_ (.A(_0773_),
    .B(_0812_),
    .Y(_0813_));
 sky130_fd_sc_hd__a21oi_1 _1188_ (.A1(_0793_),
    .A2(_0798_),
    .B1(_0811_),
    .Y(_0814_));
 sky130_fd_sc_hd__mux2_1 _1189_ (.A0(\register_file.write_data[18] ),
    .A1(\id_ex_rs1_data[18] ),
    .S(_0618_),
    .X(_0815_));
 sky130_fd_sc_hd__mux2_1 _1190_ (.A0(net380),
    .A1(_0815_),
    .S(_0620_),
    .X(_0816_));
 sky130_fd_sc_hd__o21a_1 _1191_ (.A1(_0813_),
    .A2(_0814_),
    .B1(_0816_),
    .X(_0817_));
 sky130_fd_sc_hd__nor3_1 _1192_ (.A(_0813_),
    .B(_0814_),
    .C(_0816_),
    .Y(_0818_));
 sky130_fd_sc_hd__or2_2 _1193_ (.A(_0817_),
    .B(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__o21a_1 _1194_ (.A1(_0780_),
    .A2(_0804_),
    .B1(_0805_),
    .X(_0820_));
 sky130_fd_sc_hd__o31a_1 _1195_ (.A1(_0782_),
    .A2(_0790_),
    .A3(_0806_),
    .B1(_0820_),
    .X(_0821_));
 sky130_fd_sc_hd__o21ai_1 _1196_ (.A1(_0819_),
    .A2(_0821_),
    .B1(_0592_),
    .Y(_0822_));
 sky130_fd_sc_hd__a21oi_1 _1197_ (.A1(_0819_),
    .A2(_0821_),
    .B1(_0822_),
    .Y(_0051_));
 sky130_fd_sc_hd__mux2_1 _1198_ (.A0(\register_file.write_data[19] ),
    .A1(\id_ex_rs2_data[19] ),
    .S(_0609_),
    .X(_0823_));
 sky130_fd_sc_hd__or2_1 _1199_ (.A(\dmem.address[19] ),
    .B(_0611_),
    .X(_0824_));
 sky130_fd_sc_hd__o211a_1 _1200_ (.A1(_0794_),
    .A2(_0823_),
    .B1(_0824_),
    .C1(_0613_),
    .X(_0825_));
 sky130_fd_sc_hd__xor2_2 _1201_ (.A(_0813_),
    .B(_0825_),
    .X(_0826_));
 sky130_fd_sc_hd__mux2_1 _1202_ (.A0(\register_file.write_data[19] ),
    .A1(\id_ex_rs1_data[19] ),
    .S(_0690_),
    .X(_0827_));
 sky130_fd_sc_hd__mux2_1 _1203_ (.A0(net370),
    .A1(_0827_),
    .S(_0692_),
    .X(_0828_));
 sky130_fd_sc_hd__xnor2_2 _1204_ (.A(_0826_),
    .B(_0828_),
    .Y(_0829_));
 sky130_fd_sc_hd__o21ba_1 _1205_ (.A1(_0819_),
    .A2(_0821_),
    .B1_N(_0817_),
    .X(_0830_));
 sky130_fd_sc_hd__a21oi_1 _1206_ (.A1(_0829_),
    .A2(_0830_),
    .B1(_0564_),
    .Y(_0831_));
 sky130_fd_sc_hd__o21a_1 _1207_ (.A1(_0829_),
    .A2(_0830_),
    .B1(_0831_),
    .X(_0052_));
 sky130_fd_sc_hd__or2_2 _1208_ (.A(_0812_),
    .B(_0825_),
    .X(_0832_));
 sky130_fd_sc_hd__buf_4 _1209_ (.A(_0609_),
    .X(_0833_));
 sky130_fd_sc_hd__mux2_1 _1210_ (.A0(\register_file.write_data[20] ),
    .A1(\id_ex_rs2_data[20] ),
    .S(_0833_),
    .X(_0834_));
 sky130_fd_sc_hd__buf_2 _1211_ (.A(_0611_),
    .X(_0835_));
 sky130_fd_sc_hd__or2_1 _1212_ (.A(\dmem.address[20] ),
    .B(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__clkbuf_4 _1213_ (.A(_0613_),
    .X(_0837_));
 sky130_fd_sc_hd__o211a_1 _1214_ (.A1(_0794_),
    .A2(_0834_),
    .B1(_0836_),
    .C1(_0837_),
    .X(_0838_));
 sky130_fd_sc_hd__or3_1 _1215_ (.A(_0773_),
    .B(_0832_),
    .C(_0838_),
    .X(_0839_));
 sky130_fd_sc_hd__o21ai_1 _1216_ (.A1(_0773_),
    .A2(_0832_),
    .B1(_0838_),
    .Y(_0840_));
 sky130_fd_sc_hd__or2_1 _1217_ (.A(\register_file.write_data[20] ),
    .B(_0528_),
    .X(_0841_));
 sky130_fd_sc_hd__o211a_1 _1218_ (.A1(\id_ex_rs1_data[20] ),
    .A2(_0558_),
    .B1(_0841_),
    .C1(_0532_),
    .X(_0279_));
 sky130_fd_sc_hd__a21oi_1 _1219_ (.A1(net335),
    .A2(_0556_),
    .B1(_0279_),
    .Y(_0280_));
 sky130_fd_sc_hd__a21oi_1 _1220_ (.A1(_0839_),
    .A2(_0840_),
    .B1(_0280_),
    .Y(_0281_));
 sky130_fd_sc_hd__and3_1 _1221_ (.A(_0839_),
    .B(_0840_),
    .C(_0280_),
    .X(_0282_));
 sky130_fd_sc_hd__or2_1 _1222_ (.A(_0281_),
    .B(_0282_),
    .X(_0283_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1223_ (.A(_0283_),
    .X(_0284_));
 sky130_fd_sc_hd__or4_1 _1224_ (.A(_0782_),
    .B(_0806_),
    .C(_0819_),
    .D(_0829_),
    .X(_0285_));
 sky130_fd_sc_hd__a21oi_1 _1225_ (.A1(_0826_),
    .A2(_0828_),
    .B1(_0817_),
    .Y(_0286_));
 sky130_fd_sc_hd__nor2_1 _1226_ (.A(_0826_),
    .B(_0828_),
    .Y(_0287_));
 sky130_fd_sc_hd__o32ai_4 _1227_ (.A1(_0819_),
    .A2(_0820_),
    .A3(_0829_),
    .B1(_0286_),
    .B2(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__o21ba_1 _1228_ (.A1(_0790_),
    .A2(_0285_),
    .B1_N(_0288_),
    .X(_0289_));
 sky130_fd_sc_hd__o21ai_1 _1229_ (.A1(_0284_),
    .A2(_0289_),
    .B1(_0519_),
    .Y(_0290_));
 sky130_fd_sc_hd__a21oi_1 _1230_ (.A1(_0284_),
    .A2(_0289_),
    .B1(_0290_),
    .Y(_0053_));
 sky130_fd_sc_hd__mux2_1 _1231_ (.A0(\register_file.write_data[21] ),
    .A1(\id_ex_rs2_data[21] ),
    .S(_0833_),
    .X(_0291_));
 sky130_fd_sc_hd__or2_1 _1232_ (.A(\dmem.address[21] ),
    .B(_0835_),
    .X(_0292_));
 sky130_fd_sc_hd__o211a_1 _1233_ (.A1(_0794_),
    .A2(_0291_),
    .B1(_0292_),
    .C1(_0837_),
    .X(_0293_));
 sky130_fd_sc_hd__nor2_1 _1234_ (.A(_0838_),
    .B(_0293_),
    .Y(_0294_));
 sky130_fd_sc_hd__nor3b_2 _1235_ (.A(_0773_),
    .B(_0832_),
    .C_N(_0294_),
    .Y(_0295_));
 sky130_fd_sc_hd__o31a_1 _1236_ (.A1(_0773_),
    .A2(_0832_),
    .A3(_0838_),
    .B1(_0293_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _1237_ (.A0(\register_file.write_data[21] ),
    .A1(\id_ex_rs1_data[21] ),
    .S(_0618_),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _1238_ (.A0(net322),
    .A1(_0297_),
    .S(_0620_),
    .X(_0298_));
 sky130_fd_sc_hd__o21a_1 _1239_ (.A1(_0295_),
    .A2(_0296_),
    .B1(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__or3_1 _1240_ (.A(_0295_),
    .B(_0296_),
    .C(_0298_),
    .X(_0300_));
 sky130_fd_sc_hd__nand2b_1 _1241_ (.A_N(_0299_),
    .B(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__o21ba_1 _1242_ (.A1(_0284_),
    .A2(_0289_),
    .B1_N(_0281_),
    .X(_0302_));
 sky130_fd_sc_hd__xnor2_1 _1243_ (.A(_0301_),
    .B(_0302_),
    .Y(_0303_));
 sky130_fd_sc_hd__nor2_1 _1244_ (.A(_0522_),
    .B(_0303_),
    .Y(_0054_));
 sky130_fd_sc_hd__mux2_1 _1245_ (.A0(\register_file.write_data[22] ),
    .A1(\id_ex_rs2_data[22] ),
    .S(_0833_),
    .X(_0304_));
 sky130_fd_sc_hd__or2_1 _1246_ (.A(\dmem.address[22] ),
    .B(_0835_),
    .X(_0305_));
 sky130_fd_sc_hd__o211a_1 _1247_ (.A1(_0794_),
    .A2(_0304_),
    .B1(_0305_),
    .C1(_0837_),
    .X(_0306_));
 sky130_fd_sc_hd__xor2_2 _1248_ (.A(_0295_),
    .B(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _1249_ (.A0(\register_file.write_data[22] ),
    .A1(\id_ex_rs1_data[22] ),
    .S(_0690_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _1250_ (.A0(net326),
    .A1(_0308_),
    .S(_0692_),
    .X(_0309_));
 sky130_fd_sc_hd__nand2_1 _1251_ (.A(_0307_),
    .B(_0309_),
    .Y(_0310_));
 sky130_fd_sc_hd__or2_1 _1252_ (.A(_0307_),
    .B(_0309_),
    .X(_0311_));
 sky130_fd_sc_hd__and2_1 _1253_ (.A(_0310_),
    .B(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__a21o_1 _1254_ (.A1(_0281_),
    .A2(_0300_),
    .B1(_0299_),
    .X(_0313_));
 sky130_fd_sc_hd__nor3_1 _1255_ (.A(_0284_),
    .B(_0289_),
    .C(_0301_),
    .Y(_0314_));
 sky130_fd_sc_hd__or3_1 _1256_ (.A(_0312_),
    .B(_0313_),
    .C(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__o21ai_1 _1257_ (.A1(_0313_),
    .A2(_0314_),
    .B1(_0312_),
    .Y(_0316_));
 sky130_fd_sc_hd__and3_1 _1258_ (.A(_0628_),
    .B(_0315_),
    .C(_0316_),
    .X(_0055_));
 sky130_fd_sc_hd__or4b_2 _1259_ (.A(_0773_),
    .B(_0832_),
    .C(_0306_),
    .D_N(_0294_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _1260_ (.A0(\register_file.write_data[23] ),
    .A1(\id_ex_rs2_data[23] ),
    .S(_0833_),
    .X(_0318_));
 sky130_fd_sc_hd__or2_1 _1261_ (.A(\dmem.address[23] ),
    .B(_0835_),
    .X(_0319_));
 sky130_fd_sc_hd__o211a_1 _1262_ (.A1(_0794_),
    .A2(_0318_),
    .B1(_0319_),
    .C1(_0837_),
    .X(_0320_));
 sky130_fd_sc_hd__xnor2_2 _1263_ (.A(_0317_),
    .B(_0320_),
    .Y(_0321_));
 sky130_fd_sc_hd__mux2_1 _1264_ (.A0(\register_file.write_data[23] ),
    .A1(\id_ex_rs1_data[23] ),
    .S(_0690_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _1265_ (.A0(net328),
    .A1(_0322_),
    .S(_0692_),
    .X(_0323_));
 sky130_fd_sc_hd__xnor2_2 _1266_ (.A(_0321_),
    .B(_0323_),
    .Y(_0324_));
 sky130_fd_sc_hd__a21oi_1 _1267_ (.A1(_0310_),
    .A2(_0316_),
    .B1(_0324_),
    .Y(_0325_));
 sky130_fd_sc_hd__a31o_1 _1268_ (.A1(_0310_),
    .A2(_0316_),
    .A3(_0324_),
    .B1(_0607_),
    .X(_0326_));
 sky130_fd_sc_hd__nor2_1 _1269_ (.A(_0325_),
    .B(_0326_),
    .Y(_0056_));
 sky130_fd_sc_hd__xnor2_1 _1270_ (.A(_0307_),
    .B(_0309_),
    .Y(_0327_));
 sky130_fd_sc_hd__or4_1 _1271_ (.A(_0284_),
    .B(_0301_),
    .C(_0327_),
    .D(_0324_),
    .X(_0328_));
 sky130_fd_sc_hd__a211o_1 _1272_ (.A1(_0784_),
    .A2(_0789_),
    .B1(_0285_),
    .C1(_0328_),
    .X(_0329_));
 sky130_fd_sc_hd__nor2_1 _1273_ (.A(_0327_),
    .B(_0324_),
    .Y(_0330_));
 sky130_fd_sc_hd__nor4_1 _1274_ (.A(_0284_),
    .B(_0301_),
    .C(_0327_),
    .D(_0324_),
    .Y(_0331_));
 sky130_fd_sc_hd__a22o_1 _1275_ (.A1(_0307_),
    .A2(_0309_),
    .B1(_0321_),
    .B2(_0323_),
    .X(_0332_));
 sky130_fd_sc_hd__o21a_1 _1276_ (.A1(_0321_),
    .A2(_0323_),
    .B1(_0332_),
    .X(_0333_));
 sky130_fd_sc_hd__a221oi_2 _1277_ (.A1(_0313_),
    .A2(_0330_),
    .B1(_0331_),
    .B2(_0288_),
    .C1(_0333_),
    .Y(_0334_));
 sky130_fd_sc_hd__nor2_1 _1278_ (.A(_0317_),
    .B(_0320_),
    .Y(_0335_));
 sky130_fd_sc_hd__mux2_1 _1279_ (.A0(\register_file.write_data[24] ),
    .A1(\id_ex_rs2_data[24] ),
    .S(_0833_),
    .X(_0336_));
 sky130_fd_sc_hd__or2_1 _1280_ (.A(\dmem.address[24] ),
    .B(_0835_),
    .X(_0337_));
 sky130_fd_sc_hd__o211a_1 _1281_ (.A1(_0794_),
    .A2(_0336_),
    .B1(_0337_),
    .C1(_0837_),
    .X(_0338_));
 sky130_fd_sc_hd__xnor2_1 _1282_ (.A(_0335_),
    .B(_0338_),
    .Y(_0339_));
 sky130_fd_sc_hd__mux2_1 _1283_ (.A0(\register_file.write_data[24] ),
    .A1(\id_ex_rs1_data[24] ),
    .S(_0690_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _1284_ (.A0(net430),
    .A1(_0340_),
    .S(_0692_),
    .X(_0341_));
 sky130_fd_sc_hd__xor2_1 _1285_ (.A(_0339_),
    .B(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__a31o_1 _1286_ (.A1(_0329_),
    .A2(_0334_),
    .A3(_0342_),
    .B1(_0521_),
    .X(_0343_));
 sky130_fd_sc_hd__a21o_1 _1287_ (.A1(_0329_),
    .A2(_0334_),
    .B1(_0342_),
    .X(_0344_));
 sky130_fd_sc_hd__nor2b_1 _1288_ (.A(_0343_),
    .B_N(_0344_),
    .Y(_0057_));
 sky130_fd_sc_hd__or2b_1 _1289_ (.A(_0339_),
    .B_N(_0341_),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _1290_ (.A0(\register_file.write_data[25] ),
    .A1(\id_ex_rs2_data[25] ),
    .S(_0833_),
    .X(_0346_));
 sky130_fd_sc_hd__or2_1 _1291_ (.A(\dmem.address[25] ),
    .B(_0835_),
    .X(_0347_));
 sky130_fd_sc_hd__o211a_1 _1292_ (.A1(_0794_),
    .A2(_0346_),
    .B1(_0347_),
    .C1(_0837_),
    .X(_0348_));
 sky130_fd_sc_hd__or4_1 _1293_ (.A(_0317_),
    .B(_0320_),
    .C(_0338_),
    .D(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1294_ (.A(_0349_),
    .X(_0350_));
 sky130_fd_sc_hd__o31ai_1 _1295_ (.A1(_0317_),
    .A2(_0320_),
    .A3(_0338_),
    .B1(_0348_),
    .Y(_0351_));
 sky130_fd_sc_hd__nand2_1 _1296_ (.A(_0350_),
    .B(_0351_),
    .Y(_0352_));
 sky130_fd_sc_hd__mux2_1 _1297_ (.A0(\register_file.write_data[25] ),
    .A1(\id_ex_rs1_data[25] ),
    .S(_0690_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _1298_ (.A0(net421),
    .A1(_0353_),
    .S(_0692_),
    .X(_0354_));
 sky130_fd_sc_hd__and2_1 _1299_ (.A(_0352_),
    .B(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__or2_1 _1300_ (.A(_0352_),
    .B(_0354_),
    .X(_0356_));
 sky130_fd_sc_hd__or2b_1 _1301_ (.A(_0355_),
    .B_N(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__a21oi_1 _1302_ (.A1(_0345_),
    .A2(_0344_),
    .B1(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__a31o_1 _1303_ (.A1(_0345_),
    .A2(_0344_),
    .A3(_0357_),
    .B1(_0607_),
    .X(_0359_));
 sky130_fd_sc_hd__nor2_1 _1304_ (.A(_0358_),
    .B(_0359_),
    .Y(_0058_));
 sky130_fd_sc_hd__a211o_1 _1305_ (.A1(_0329_),
    .A2(_0334_),
    .B1(_0342_),
    .C1(_0357_),
    .X(_0360_));
 sky130_fd_sc_hd__and2b_1 _1306_ (.A_N(_0345_),
    .B(_0356_),
    .X(_0361_));
 sky130_fd_sc_hd__nor2_1 _1307_ (.A(_0355_),
    .B(_0361_),
    .Y(_0362_));
 sky130_fd_sc_hd__mux2_1 _1308_ (.A0(\register_file.write_data[26] ),
    .A1(\id_ex_rs2_data[26] ),
    .S(_0833_),
    .X(_0363_));
 sky130_fd_sc_hd__or2_1 _1309_ (.A(net324),
    .B(_0835_),
    .X(_0364_));
 sky130_fd_sc_hd__o211a_1 _1310_ (.A1(_0794_),
    .A2(_0363_),
    .B1(_0364_),
    .C1(_0837_),
    .X(_0365_));
 sky130_fd_sc_hd__xnor2_1 _1311_ (.A(_0350_),
    .B(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__mux2_1 _1312_ (.A0(net410),
    .A1(net495),
    .S(_0690_),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _1313_ (.A0(net324),
    .A1(_0367_),
    .S(_0692_),
    .X(_0368_));
 sky130_fd_sc_hd__and2_1 _1314_ (.A(_0366_),
    .B(_0368_),
    .X(_0369_));
 sky130_fd_sc_hd__or2_1 _1315_ (.A(_0366_),
    .B(_0368_),
    .X(_0370_));
 sky130_fd_sc_hd__or2b_1 _1316_ (.A(_0369_),
    .B_N(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__a21oi_1 _1317_ (.A1(_0360_),
    .A2(_0362_),
    .B1(_0371_),
    .Y(_0372_));
 sky130_fd_sc_hd__a31o_1 _1318_ (.A1(_0371_),
    .A2(_0360_),
    .A3(_0362_),
    .B1(_0607_),
    .X(_0373_));
 sky130_fd_sc_hd__nor2_1 _1319_ (.A(_0372_),
    .B(_0373_),
    .Y(_0059_));
 sky130_fd_sc_hd__mux2_1 _1320_ (.A0(\register_file.write_data[27] ),
    .A1(\id_ex_rs2_data[27] ),
    .S(_0833_),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_1 _1321_ (.A0(net200),
    .A1(_0374_),
    .S(_0835_),
    .X(_0375_));
 sky130_fd_sc_hd__nand2_1 _1322_ (.A(_0837_),
    .B(_0375_),
    .Y(_0376_));
 sky130_fd_sc_hd__inv_2 _1323_ (.A(_0376_),
    .Y(_0377_));
 sky130_fd_sc_hd__or3_1 _1324_ (.A(_0350_),
    .B(_0365_),
    .C(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__o21ai_1 _1325_ (.A1(_0350_),
    .A2(_0365_),
    .B1(_0377_),
    .Y(_0379_));
 sky130_fd_sc_hd__mux2_1 _1326_ (.A0(\register_file.write_data[27] ),
    .A1(\id_ex_rs1_data[27] ),
    .S(_0690_),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_1 _1327_ (.A0(net200),
    .A1(_0380_),
    .S(_0692_),
    .X(_0381_));
 sky130_fd_sc_hd__inv_2 _1328_ (.A(_0381_),
    .Y(_0382_));
 sky130_fd_sc_hd__a21oi_1 _1329_ (.A1(_0378_),
    .A2(_0379_),
    .B1(_0382_),
    .Y(_0383_));
 sky130_fd_sc_hd__nand3_1 _1330_ (.A(_0378_),
    .B(_0379_),
    .C(_0382_),
    .Y(_0384_));
 sky130_fd_sc_hd__and2b_1 _1331_ (.A_N(_0383_),
    .B(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__or2_1 _1332_ (.A(_0369_),
    .B(_0372_),
    .X(_0386_));
 sky130_fd_sc_hd__a21oi_1 _1333_ (.A1(_0385_),
    .A2(_0386_),
    .B1(_0564_),
    .Y(_0387_));
 sky130_fd_sc_hd__o21a_1 _1334_ (.A1(_0385_),
    .A2(_0386_),
    .B1(_0387_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _1335_ (.A0(\register_file.write_data[28] ),
    .A1(\id_ex_rs2_data[28] ),
    .S(_0833_),
    .X(_0388_));
 sky130_fd_sc_hd__or2_1 _1336_ (.A(\dmem.address[28] ),
    .B(_0835_),
    .X(_0389_));
 sky130_fd_sc_hd__o211a_1 _1337_ (.A1(_0794_),
    .A2(_0388_),
    .B1(_0389_),
    .C1(_0837_),
    .X(_0390_));
 sky130_fd_sc_hd__xnor2_1 _1338_ (.A(_0378_),
    .B(_0390_),
    .Y(_0391_));
 sky130_fd_sc_hd__mux2_1 _1339_ (.A0(net351),
    .A1(\id_ex_rs1_data[28] ),
    .S(_0690_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _1340_ (.A0(net435),
    .A1(_0392_),
    .S(_0692_),
    .X(_0393_));
 sky130_fd_sc_hd__xnor2_1 _1341_ (.A(_0391_),
    .B(_0393_),
    .Y(_0394_));
 sky130_fd_sc_hd__a21oi_1 _1342_ (.A1(_0369_),
    .A2(_0384_),
    .B1(_0383_),
    .Y(_0395_));
 sky130_fd_sc_hd__a21oi_1 _1343_ (.A1(_0370_),
    .A2(_0384_),
    .B1(_0383_),
    .Y(_0396_));
 sky130_fd_sc_hd__a31o_1 _1344_ (.A1(_0360_),
    .A2(_0362_),
    .A3(_0395_),
    .B1(_0396_),
    .X(_0397_));
 sky130_fd_sc_hd__nor2_1 _1345_ (.A(_0394_),
    .B(_0397_),
    .Y(_0398_));
 sky130_fd_sc_hd__or2_1 _1346_ (.A(_0521_),
    .B(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__a21oi_1 _1347_ (.A1(_0394_),
    .A2(_0397_),
    .B1(_0399_),
    .Y(_0061_));
 sky130_fd_sc_hd__and2_1 _1348_ (.A(_0391_),
    .B(_0393_),
    .X(_0400_));
 sky130_fd_sc_hd__or4_1 _1349_ (.A(_0350_),
    .B(_0365_),
    .C(_0377_),
    .D(_0390_),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_1 _1350_ (.A0(\register_file.write_data[29] ),
    .A1(\id_ex_rs2_data[29] ),
    .S(_0833_),
    .X(_0402_));
 sky130_fd_sc_hd__or2_1 _1351_ (.A(\dmem.address[29] ),
    .B(_0835_),
    .X(_0403_));
 sky130_fd_sc_hd__o211a_1 _1352_ (.A1(_0794_),
    .A2(_0402_),
    .B1(_0403_),
    .C1(_0837_),
    .X(_0404_));
 sky130_fd_sc_hd__xnor2_1 _1353_ (.A(_0401_),
    .B(_0404_),
    .Y(_0405_));
 sky130_fd_sc_hd__mux2_1 _1354_ (.A0(net536),
    .A1(\id_ex_rs1_data[29] ),
    .S(_0690_),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_1 _1355_ (.A0(net437),
    .A1(_0406_),
    .S(_0692_),
    .X(_0407_));
 sky130_fd_sc_hd__xnor2_1 _1356_ (.A(_0405_),
    .B(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__nor3b_1 _1357_ (.A(_0400_),
    .B(_0398_),
    .C_N(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__o21ba_1 _1358_ (.A1(_0400_),
    .A2(_0398_),
    .B1_N(_0408_),
    .X(_0410_));
 sky130_fd_sc_hd__nor3_1 _1359_ (.A(_0522_),
    .B(_0409_),
    .C(_0410_),
    .Y(_0062_));
 sky130_fd_sc_hd__buf_1 _1360_ (.A(_0519_),
    .X(_0411_));
 sky130_fd_sc_hd__nand2_1 _1361_ (.A(_0405_),
    .B(_0407_),
    .Y(_0412_));
 sky130_fd_sc_hd__nor2_1 _1362_ (.A(_0401_),
    .B(_0404_),
    .Y(_0413_));
 sky130_fd_sc_hd__mux2_1 _1363_ (.A0(\register_file.write_data[30] ),
    .A1(\id_ex_rs2_data[30] ),
    .S(_0833_),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _1364_ (.A0(net418),
    .A1(_0414_),
    .S(_0835_),
    .X(_0415_));
 sky130_fd_sc_hd__nand2_1 _1365_ (.A(_0837_),
    .B(_0415_),
    .Y(_0416_));
 sky130_fd_sc_hd__xor2_1 _1366_ (.A(_0413_),
    .B(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _1367_ (.A0(\register_file.write_data[30] ),
    .A1(\id_ex_rs1_data[30] ),
    .S(_0690_),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _1368_ (.A0(net418),
    .A1(_0418_),
    .S(_0692_),
    .X(_0419_));
 sky130_fd_sc_hd__or2b_1 _1369_ (.A(_0417_),
    .B_N(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__or2b_1 _1370_ (.A(_0419_),
    .B_N(_0417_),
    .X(_0421_));
 sky130_fd_sc_hd__nand2_1 _1371_ (.A(_0420_),
    .B(_0421_),
    .Y(_0422_));
 sky130_fd_sc_hd__or2_1 _1372_ (.A(_0394_),
    .B(_0408_),
    .X(_0423_));
 sky130_fd_sc_hd__a311o_1 _1373_ (.A1(_0360_),
    .A2(_0362_),
    .A3(_0395_),
    .B1(_0396_),
    .C1(_0423_),
    .X(_0424_));
 sky130_fd_sc_hd__o21ai_1 _1374_ (.A1(_0405_),
    .A2(_0407_),
    .B1(_0400_),
    .Y(_0425_));
 sky130_fd_sc_hd__nand4_1 _1375_ (.A(_0412_),
    .B(_0422_),
    .C(_0424_),
    .D(_0425_),
    .Y(_0426_));
 sky130_fd_sc_hd__a31o_1 _1376_ (.A1(_0412_),
    .A2(_0424_),
    .A3(_0425_),
    .B1(_0422_),
    .X(_0427_));
 sky130_fd_sc_hd__and3_1 _1377_ (.A(_0411_),
    .B(_0426_),
    .C(_0427_),
    .X(_0063_));
 sky130_fd_sc_hd__nand2_1 _1378_ (.A(_0413_),
    .B(_0416_),
    .Y(_0428_));
 sky130_fd_sc_hd__mux2_1 _1379_ (.A0(\register_file.write_data[31] ),
    .A1(\id_ex_rs2_data[31] ),
    .S(_0833_),
    .X(_0429_));
 sky130_fd_sc_hd__or2_1 _1380_ (.A(net429),
    .B(_0835_),
    .X(_0430_));
 sky130_fd_sc_hd__o211a_1 _1381_ (.A1(_0794_),
    .A2(_0429_),
    .B1(_0430_),
    .C1(_0837_),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _1382_ (.A0(\register_file.write_data[31] ),
    .A1(\id_ex_rs1_data[31] ),
    .S(_0690_),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_1 _1383_ (.A0(net429),
    .A1(_0432_),
    .S(_0692_),
    .X(_0433_));
 sky130_fd_sc_hd__xnor2_1 _1384_ (.A(_0431_),
    .B(_0433_),
    .Y(_0434_));
 sky130_fd_sc_hd__xnor2_1 _1385_ (.A(_0428_),
    .B(_0434_),
    .Y(_0435_));
 sky130_fd_sc_hd__a21oi_1 _1386_ (.A1(_0420_),
    .A2(_0427_),
    .B1(_0435_),
    .Y(_0436_));
 sky130_fd_sc_hd__a31o_1 _1387_ (.A1(_0420_),
    .A2(_0427_),
    .A3(_0435_),
    .B1(_0607_),
    .X(_0437_));
 sky130_fd_sc_hd__nor2_1 _1388_ (.A(_0436_),
    .B(_0437_),
    .Y(_0064_));
 sky130_fd_sc_hd__and2_1 _1389_ (.A(_0525_),
    .B(net412),
    .X(_0065_));
 sky130_fd_sc_hd__and2_1 _1390_ (.A(_0525_),
    .B(net413),
    .X(_0066_));
 sky130_fd_sc_hd__and2_1 _1391_ (.A(net533),
    .B(_0628_),
    .X(_0067_));
 sky130_fd_sc_hd__and2_1 _1392_ (.A(net459),
    .B(_0628_),
    .X(_0068_));
 sky130_fd_sc_hd__or3_1 _1393_ (.A(net105),
    .B(net134),
    .C(net106),
    .X(_0438_));
 sky130_fd_sc_hd__or4_1 _1394_ (.A(net131),
    .B(net130),
    .C(net471),
    .D(net132),
    .X(_0439_));
 sky130_fd_sc_hd__or4_4 _1395_ (.A(reset),
    .B(net129),
    .C(net499),
    .D(net472),
    .X(_0440_));
 sky130_fd_sc_hd__nor3b_1 _1396_ (.A(_0440_),
    .B(net330),
    .C_N(net434),
    .Y(_0069_));
 sky130_fd_sc_hd__buf_2 _1397_ (.A(net337),
    .X(_0441_));
 sky130_fd_sc_hd__and2_1 _1398_ (.A(_0441_),
    .B(_0628_),
    .X(_0070_));
 sky130_fd_sc_hd__and2_1 _1399_ (.A(_0519_),
    .B(net490),
    .X(_0071_));
 sky130_fd_sc_hd__and2_1 _1400_ (.A(_0525_),
    .B(net408),
    .X(_0072_));
 sky130_fd_sc_hd__and2_1 _1401_ (.A(_0525_),
    .B(net404),
    .X(_0073_));
 sky130_fd_sc_hd__and2_1 _1402_ (.A(_0525_),
    .B(net534),
    .X(_0074_));
 sky130_fd_sc_hd__buf_1 _1403_ (.A(_0519_),
    .X(_0442_));
 sky130_fd_sc_hd__and2_1 _1404_ (.A(_0442_),
    .B(net431),
    .X(_0075_));
 sky130_fd_sc_hd__and2_1 _1405_ (.A(_0442_),
    .B(net333),
    .X(_0076_));
 sky130_fd_sc_hd__and2_1 _1406_ (.A(net441),
    .B(_0628_),
    .X(_0077_));
 sky130_fd_sc_hd__and2_1 _1407_ (.A(net433),
    .B(_0628_),
    .X(_0078_));
 sky130_fd_sc_hd__nor2_1 _1408_ (.A(_0522_),
    .B(net434),
    .Y(_0079_));
 sky130_fd_sc_hd__xnor2_1 _1409_ (.A(net330),
    .B(net434),
    .Y(_0443_));
 sky130_fd_sc_hd__nor2_1 _1410_ (.A(_0522_),
    .B(_0443_),
    .Y(_0080_));
 sky130_fd_sc_hd__a21oi_1 _1411_ (.A1(net330),
    .A2(net125),
    .B1(net129),
    .Y(_0444_));
 sky130_fd_sc_hd__a31o_1 _1412_ (.A1(net129),
    .A2(net330),
    .A3(net125),
    .B1(_0521_),
    .X(_0445_));
 sky130_fd_sc_hd__nor2_1 _1413_ (.A(net331),
    .B(_0445_),
    .Y(_0081_));
 sky130_fd_sc_hd__and4_1 _1414_ (.A(net525),
    .B(net401),
    .C(net330),
    .D(net125),
    .X(_0446_));
 sky130_fd_sc_hd__a31o_1 _1415_ (.A1(net129),
    .A2(net330),
    .A3(net125),
    .B1(net401),
    .X(_0447_));
 sky130_fd_sc_hd__nand2_1 _1416_ (.A(_0592_),
    .B(net402),
    .Y(_0448_));
 sky130_fd_sc_hd__nor2_1 _1417_ (.A(_0446_),
    .B(_0448_),
    .Y(_0082_));
 sky130_fd_sc_hd__a21oi_1 _1418_ (.A1(net500),
    .A2(_0446_),
    .B1(_0564_),
    .Y(_0449_));
 sky130_fd_sc_hd__o21a_1 _1419_ (.A1(net500),
    .A2(_0446_),
    .B1(_0449_),
    .X(_0083_));
 sky130_fd_sc_hd__a21oi_1 _1420_ (.A1(net500),
    .A2(_0446_),
    .B1(net491),
    .Y(_0450_));
 sky130_fd_sc_hd__and3_1 _1421_ (.A(net131),
    .B(net491),
    .C(_0446_),
    .X(_0451_));
 sky130_fd_sc_hd__nor3_1 _1422_ (.A(_0522_),
    .B(_0450_),
    .C(net492),
    .Y(_0084_));
 sky130_fd_sc_hd__buf_1 _1423_ (.A(_0521_),
    .X(_0452_));
 sky130_fd_sc_hd__and4_1 _1424_ (.A(net500),
    .B(net471),
    .C(net491),
    .D(_0446_),
    .X(_0453_));
 sky130_fd_sc_hd__nor2_1 _1425_ (.A(_0452_),
    .B(_0453_),
    .Y(_0454_));
 sky130_fd_sc_hd__o21a_1 _1426_ (.A1(net471),
    .A2(net492),
    .B1(_0454_),
    .X(_0085_));
 sky130_fd_sc_hd__a21oi_1 _1427_ (.A1(net505),
    .A2(_0453_),
    .B1(_0564_),
    .Y(_0455_));
 sky130_fd_sc_hd__o21a_1 _1428_ (.A1(net505),
    .A2(_0453_),
    .B1(_0455_),
    .X(_0086_));
 sky130_fd_sc_hd__a21oi_1 _1429_ (.A1(net134),
    .A2(_0453_),
    .B1(net502),
    .Y(_0456_));
 sky130_fd_sc_hd__and3_1 _1430_ (.A(net502),
    .B(net505),
    .C(_0453_),
    .X(_0457_));
 sky130_fd_sc_hd__nor3_1 _1431_ (.A(_0522_),
    .B(net503),
    .C(_0457_),
    .Y(_0087_));
 sky130_fd_sc_hd__and4_1 _1432_ (.A(net502),
    .B(net505),
    .C(net498),
    .D(_0453_),
    .X(_0458_));
 sky130_fd_sc_hd__nor2_1 _1433_ (.A(_0452_),
    .B(_0458_),
    .Y(_0459_));
 sky130_fd_sc_hd__o21a_1 _1434_ (.A1(net498),
    .A2(_0457_),
    .B1(_0459_),
    .X(_0088_));
 sky130_fd_sc_hd__a21oi_1 _1435_ (.A1(net457),
    .A2(_0458_),
    .B1(_0564_),
    .Y(_0460_));
 sky130_fd_sc_hd__o21a_1 _1436_ (.A1(net457),
    .A2(_0458_),
    .B1(_0460_),
    .X(_0089_));
 sky130_fd_sc_hd__a21oi_1 _1437_ (.A1(net457),
    .A2(_0458_),
    .B1(net415),
    .Y(_0461_));
 sky130_fd_sc_hd__and3_1 _1438_ (.A(net107),
    .B(net415),
    .C(_0458_),
    .X(_0462_));
 sky130_fd_sc_hd__nor3_1 _1439_ (.A(_0522_),
    .B(net458),
    .C(net416),
    .Y(_0090_));
 sky130_fd_sc_hd__and2_1 _1440_ (.A(net109),
    .B(net416),
    .X(_0463_));
 sky130_fd_sc_hd__nor2_1 _1441_ (.A(_0452_),
    .B(_0463_),
    .Y(_0464_));
 sky130_fd_sc_hd__o21a_1 _1442_ (.A1(net109),
    .A2(net416),
    .B1(_0464_),
    .X(_0091_));
 sky130_fd_sc_hd__a21oi_1 _1443_ (.A1(net514),
    .A2(_0463_),
    .B1(_0564_),
    .Y(_0465_));
 sky130_fd_sc_hd__o21a_1 _1444_ (.A1(net514),
    .A2(_0463_),
    .B1(_0465_),
    .X(_0092_));
 sky130_fd_sc_hd__a21oi_1 _1445_ (.A1(net110),
    .A2(_0463_),
    .B1(net466),
    .Y(_0466_));
 sky130_fd_sc_hd__and3_1 _1446_ (.A(net518),
    .B(net466),
    .C(_0463_),
    .X(_0467_));
 sky130_fd_sc_hd__nor3_1 _1447_ (.A(_0522_),
    .B(net467),
    .C(_0467_),
    .Y(_0093_));
 sky130_fd_sc_hd__and2_1 _1448_ (.A(net451),
    .B(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__nor2_1 _1449_ (.A(_0452_),
    .B(_0468_),
    .Y(_0469_));
 sky130_fd_sc_hd__o21a_1 _1450_ (.A1(net451),
    .A2(_0467_),
    .B1(_0469_),
    .X(_0094_));
 sky130_fd_sc_hd__a21oi_1 _1451_ (.A1(net516),
    .A2(_0468_),
    .B1(_0564_),
    .Y(_0470_));
 sky130_fd_sc_hd__o21a_1 _1452_ (.A1(net516),
    .A2(_0468_),
    .B1(_0470_),
    .X(_0095_));
 sky130_fd_sc_hd__a21oi_1 _1453_ (.A1(net113),
    .A2(_0468_),
    .B1(net463),
    .Y(_0471_));
 sky130_fd_sc_hd__and3_1 _1454_ (.A(net113),
    .B(net463),
    .C(_0468_),
    .X(_0472_));
 sky130_fd_sc_hd__nor3_1 _1455_ (.A(_0522_),
    .B(net464),
    .C(_0472_),
    .Y(_0096_));
 sky130_fd_sc_hd__and2_1 _1456_ (.A(net447),
    .B(net517),
    .X(_0473_));
 sky130_fd_sc_hd__nor2_1 _1457_ (.A(_0452_),
    .B(_0473_),
    .Y(_0474_));
 sky130_fd_sc_hd__o21a_1 _1458_ (.A1(net447),
    .A2(_0472_),
    .B1(_0474_),
    .X(_0097_));
 sky130_fd_sc_hd__a21oi_1 _1459_ (.A1(net426),
    .A2(_0473_),
    .B1(_0452_),
    .Y(_0475_));
 sky130_fd_sc_hd__o21a_1 _1460_ (.A1(net426),
    .A2(_0473_),
    .B1(_0475_),
    .X(_0098_));
 sky130_fd_sc_hd__a21oi_1 _1461_ (.A1(net426),
    .A2(_0473_),
    .B1(net117),
    .Y(_0476_));
 sky130_fd_sc_hd__and3_1 _1462_ (.A(net426),
    .B(net117),
    .C(_0473_),
    .X(_0477_));
 sky130_fd_sc_hd__nor3_1 _1463_ (.A(_0564_),
    .B(net427),
    .C(_0477_),
    .Y(_0099_));
 sky130_fd_sc_hd__and2_1 _1464_ (.A(net449),
    .B(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__nor2_1 _1465_ (.A(_0452_),
    .B(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__o21a_1 _1466_ (.A1(net449),
    .A2(_0477_),
    .B1(_0479_),
    .X(_0100_));
 sky130_fd_sc_hd__a21oi_1 _1467_ (.A1(net512),
    .A2(_0478_),
    .B1(_0452_),
    .Y(_0480_));
 sky130_fd_sc_hd__o21a_1 _1468_ (.A1(net512),
    .A2(_0478_),
    .B1(_0480_),
    .X(_0101_));
 sky130_fd_sc_hd__a21oi_1 _1469_ (.A1(net119),
    .A2(_0478_),
    .B1(net460),
    .Y(_0481_));
 sky130_fd_sc_hd__and3_1 _1470_ (.A(net541),
    .B(net460),
    .C(_0478_),
    .X(_0482_));
 sky130_fd_sc_hd__nor3_1 _1471_ (.A(_0564_),
    .B(net461),
    .C(_0482_),
    .Y(_0102_));
 sky130_fd_sc_hd__and2_1 _1472_ (.A(net455),
    .B(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__nor2_1 _1473_ (.A(_0452_),
    .B(_0483_),
    .Y(_0484_));
 sky130_fd_sc_hd__o21a_1 _1474_ (.A1(net455),
    .A2(_0482_),
    .B1(_0484_),
    .X(_0103_));
 sky130_fd_sc_hd__a21oi_1 _1475_ (.A1(net511),
    .A2(_0483_),
    .B1(_0452_),
    .Y(_0485_));
 sky130_fd_sc_hd__o21a_1 _1476_ (.A1(net511),
    .A2(_0483_),
    .B1(_0485_),
    .X(_0104_));
 sky130_fd_sc_hd__a21oi_1 _1477_ (.A1(net122),
    .A2(_0483_),
    .B1(net474),
    .Y(_0486_));
 sky130_fd_sc_hd__and3_1 _1478_ (.A(net540),
    .B(net474),
    .C(_0483_),
    .X(_0487_));
 sky130_fd_sc_hd__nor3_1 _1479_ (.A(_0564_),
    .B(net475),
    .C(_0487_),
    .Y(_0105_));
 sky130_fd_sc_hd__and2_1 _1480_ (.A(net484),
    .B(_0487_),
    .X(_0488_));
 sky130_fd_sc_hd__nor2_1 _1481_ (.A(_0452_),
    .B(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__o21a_1 _1482_ (.A1(net484),
    .A2(_0487_),
    .B1(_0489_),
    .X(_0106_));
 sky130_fd_sc_hd__and3_1 _1483_ (.A(net484),
    .B(net479),
    .C(_0487_),
    .X(_0490_));
 sky130_fd_sc_hd__nor2_1 _1484_ (.A(_0607_),
    .B(_0490_),
    .Y(_0491_));
 sky130_fd_sc_hd__o21a_1 _1485_ (.A1(net479),
    .A2(_0488_),
    .B1(_0491_),
    .X(_0107_));
 sky130_fd_sc_hd__a21oi_1 _1486_ (.A1(net497),
    .A2(_0490_),
    .B1(_0452_),
    .Y(_0492_));
 sky130_fd_sc_hd__o21a_1 _1487_ (.A1(net497),
    .A2(_0490_),
    .B1(_0492_),
    .X(_0108_));
 sky130_fd_sc_hd__or3b_4 _1488_ (.A(_0526_),
    .B(reset),
    .C_N(mem_wb_valid),
    .X(_0493_));
 sky130_fd_sc_hd__inv_2 _1489_ (.A(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__and3_1 _1490_ (.A(net313),
    .B(net308),
    .C(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__clkbuf_4 _1491_ (.A(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__clkbuf_4 _1492_ (.A(_0496_),
    .X(_0497_));
 sky130_fd_sc_hd__nor2_4 _1493_ (.A(_0521_),
    .B(_0496_),
    .Y(_0498_));
 sky130_fd_sc_hd__clkbuf_4 _1494_ (.A(_0498_),
    .X(_0499_));
 sky130_fd_sc_hd__a22o_1 _1495_ (.A1(net300),
    .A2(_0497_),
    .B1(_0499_),
    .B2(net442),
    .X(_0109_));
 sky130_fd_sc_hd__a22o_1 _1496_ (.A1(net294),
    .A2(_0497_),
    .B1(_0499_),
    .B2(net444),
    .X(_0110_));
 sky130_fd_sc_hd__a22o_1 _1497_ (.A1(net290),
    .A2(_0497_),
    .B1(_0499_),
    .B2(net445),
    .X(_0111_));
 sky130_fd_sc_hd__a22o_1 _1498_ (.A1(net292),
    .A2(_0497_),
    .B1(_0499_),
    .B2(net443),
    .X(_0112_));
 sky130_fd_sc_hd__a22o_1 _1499_ (.A1(\register_file.write_data[4] ),
    .A2(_0497_),
    .B1(_0499_),
    .B2(net454),
    .X(_0113_));
 sky130_fd_sc_hd__a22o_1 _1500_ (.A1(\register_file.write_data[5] ),
    .A2(_0497_),
    .B1(_0499_),
    .B2(net453),
    .X(_0114_));
 sky130_fd_sc_hd__a22o_1 _1501_ (.A1(\register_file.write_data[6] ),
    .A2(_0497_),
    .B1(_0499_),
    .B2(net440),
    .X(_0115_));
 sky130_fd_sc_hd__a22o_1 _1502_ (.A1(\register_file.write_data[7] ),
    .A2(_0497_),
    .B1(_0499_),
    .B2(net446),
    .X(_0116_));
 sky130_fd_sc_hd__a22o_1 _1503_ (.A1(net296),
    .A2(_0497_),
    .B1(_0499_),
    .B2(net391),
    .X(_0117_));
 sky130_fd_sc_hd__a22o_1 _1504_ (.A1(net302),
    .A2(_0497_),
    .B1(_0499_),
    .B2(net394),
    .X(_0118_));
 sky130_fd_sc_hd__a22o_1 _1505_ (.A1(net210),
    .A2(_0497_),
    .B1(_0499_),
    .B2(net387),
    .X(_0119_));
 sky130_fd_sc_hd__a22o_1 _1506_ (.A1(net218),
    .A2(_0497_),
    .B1(_0499_),
    .B2(net388),
    .X(_0120_));
 sky130_fd_sc_hd__clkbuf_4 _1507_ (.A(_0496_),
    .X(_0500_));
 sky130_fd_sc_hd__clkbuf_4 _1508_ (.A(_0498_),
    .X(_0501_));
 sky130_fd_sc_hd__a22o_1 _1509_ (.A1(net212),
    .A2(_0500_),
    .B1(_0501_),
    .B2(net240),
    .X(_0121_));
 sky130_fd_sc_hd__a22o_1 _1510_ (.A1(net220),
    .A2(_0500_),
    .B1(_0501_),
    .B2(net246),
    .X(_0122_));
 sky130_fd_sc_hd__a22o_1 _1511_ (.A1(net208),
    .A2(_0500_),
    .B1(_0501_),
    .B2(net234),
    .X(_0123_));
 sky130_fd_sc_hd__a22o_1 _1512_ (.A1(net204),
    .A2(_0500_),
    .B1(_0501_),
    .B2(net238),
    .X(_0124_));
 sky130_fd_sc_hd__a22o_1 _1513_ (.A1(net206),
    .A2(_0500_),
    .B1(_0501_),
    .B2(net236),
    .X(_0125_));
 sky130_fd_sc_hd__a22o_1 _1514_ (.A1(net214),
    .A2(_0500_),
    .B1(_0501_),
    .B2(net242),
    .X(_0126_));
 sky130_fd_sc_hd__a22o_1 _1515_ (.A1(net216),
    .A2(_0500_),
    .B1(_0501_),
    .B2(net244),
    .X(_0127_));
 sky130_fd_sc_hd__a22o_1 _1516_ (.A1(net202),
    .A2(_0500_),
    .B1(_0501_),
    .B2(net232),
    .X(_0128_));
 sky130_fd_sc_hd__a22o_1 _1517_ (.A1(net228),
    .A2(_0500_),
    .B1(_0501_),
    .B2(net288),
    .X(_0129_));
 sky130_fd_sc_hd__a22o_1 _1518_ (.A1(net226),
    .A2(_0500_),
    .B1(_0501_),
    .B2(net286),
    .X(_0130_));
 sky130_fd_sc_hd__a22o_1 _1519_ (.A1(net224),
    .A2(_0500_),
    .B1(_0501_),
    .B2(net248),
    .X(_0131_));
 sky130_fd_sc_hd__a22o_1 _1520_ (.A1(net222),
    .A2(_0500_),
    .B1(_0501_),
    .B2(net250),
    .X(_0132_));
 sky130_fd_sc_hd__a22o_1 _1521_ (.A1(net282),
    .A2(_0496_),
    .B1(_0498_),
    .B2(net81),
    .X(_0133_));
 sky130_fd_sc_hd__a22o_1 _1522_ (.A1(net278),
    .A2(_0496_),
    .B1(_0498_),
    .B2(net82),
    .X(_0134_));
 sky130_fd_sc_hd__a22o_1 _1523_ (.A1(net280),
    .A2(_0496_),
    .B1(_0498_),
    .B2(net83),
    .X(_0135_));
 sky130_fd_sc_hd__a22o_1 _1524_ (.A1(\register_file.write_data[27] ),
    .A2(_0496_),
    .B1(_0498_),
    .B2(net469),
    .X(_0136_));
 sky130_fd_sc_hd__a22o_1 _1525_ (.A1(net351),
    .A2(_0496_),
    .B1(_0498_),
    .B2(net85),
    .X(_0137_));
 sky130_fd_sc_hd__a22o_1 _1526_ (.A1(net341),
    .A2(_0496_),
    .B1(_0498_),
    .B2(net86),
    .X(_0138_));
 sky130_fd_sc_hd__a22o_1 _1527_ (.A1(net372),
    .A2(_0496_),
    .B1(_0498_),
    .B2(net392),
    .X(_0139_));
 sky130_fd_sc_hd__a22o_1 _1528_ (.A1(net378),
    .A2(_0496_),
    .B1(_0498_),
    .B2(net393),
    .X(_0140_));
 sky130_fd_sc_hd__nor3b_2 _1529_ (.A(net100),
    .B(net404),
    .C_N(_0071_),
    .Y(_0502_));
 sky130_fd_sc_hd__clkbuf_2 _1530_ (.A(net140),
    .X(_0503_));
 sky130_fd_sc_hd__and2_1 _1531_ (.A(net33),
    .B(_0503_),
    .X(_0141_));
 sky130_fd_sc_hd__and2_1 _1532_ (.A(net44),
    .B(_0503_),
    .X(_0142_));
 sky130_fd_sc_hd__and2_1 _1533_ (.A(net419),
    .B(_0503_),
    .X(_0143_));
 sky130_fd_sc_hd__and2_1 _1534_ (.A(net58),
    .B(_0503_),
    .X(_0144_));
 sky130_fd_sc_hd__and2_1 _1535_ (.A(net389),
    .B(_0503_),
    .X(_0145_));
 sky130_fd_sc_hd__and2_1 _1536_ (.A(net488),
    .B(_0503_),
    .X(_0146_));
 sky130_fd_sc_hd__and2_1 _1537_ (.A(net366),
    .B(_0503_),
    .X(_0147_));
 sky130_fd_sc_hd__and2_1 _1538_ (.A(net368),
    .B(_0503_),
    .X(_0148_));
 sky130_fd_sc_hd__and2_1 _1539_ (.A(net537),
    .B(_0503_),
    .X(_0149_));
 sky130_fd_sc_hd__and2_1 _1540_ (.A(net383),
    .B(_0503_),
    .X(_0150_));
 sky130_fd_sc_hd__and2_1 _1541_ (.A(net270),
    .B(_0503_),
    .X(_0151_));
 sky130_fd_sc_hd__and2_1 _1542_ (.A(net276),
    .B(_0503_),
    .X(_0152_));
 sky130_fd_sc_hd__clkbuf_2 _1543_ (.A(net140),
    .X(_0504_));
 sky130_fd_sc_hd__and2_1 _1544_ (.A(net272),
    .B(_0504_),
    .X(_0153_));
 sky130_fd_sc_hd__and2_1 _1545_ (.A(net274),
    .B(_0504_),
    .X(_0154_));
 sky130_fd_sc_hd__and2_1 _1546_ (.A(net262),
    .B(_0504_),
    .X(_0155_));
 sky130_fd_sc_hd__and2_1 _1547_ (.A(net256),
    .B(_0504_),
    .X(_0156_));
 sky130_fd_sc_hd__and2_1 _1548_ (.A(net254),
    .B(_0504_),
    .X(_0157_));
 sky130_fd_sc_hd__and2_1 _1549_ (.A(net268),
    .B(_0504_),
    .X(_0158_));
 sky130_fd_sc_hd__and2_1 _1550_ (.A(net266),
    .B(_0504_),
    .X(_0159_));
 sky130_fd_sc_hd__and2_1 _1551_ (.A(net252),
    .B(_0504_),
    .X(_0160_));
 sky130_fd_sc_hd__and2_1 _1552_ (.A(net320),
    .B(_0504_),
    .X(_0161_));
 sky130_fd_sc_hd__and2_1 _1553_ (.A(net316),
    .B(_0504_),
    .X(_0162_));
 sky130_fd_sc_hd__and2_1 _1554_ (.A(net304),
    .B(_0504_),
    .X(_0163_));
 sky130_fd_sc_hd__and2_1 _1555_ (.A(net306),
    .B(_0504_),
    .X(_0164_));
 sky130_fd_sc_hd__and2_1 _1556_ (.A(net318),
    .B(net140),
    .X(_0165_));
 sky130_fd_sc_hd__and2_1 _1557_ (.A(net539),
    .B(net140),
    .X(_0166_));
 sky130_fd_sc_hd__and2_1 _1558_ (.A(net349),
    .B(net140),
    .X(_0167_));
 sky130_fd_sc_hd__and2_1 _1559_ (.A(net347),
    .B(net140),
    .X(_0168_));
 sky130_fd_sc_hd__and2_1 _1560_ (.A(net357),
    .B(net140),
    .X(_0169_));
 sky130_fd_sc_hd__and2_1 _1561_ (.A(net343),
    .B(net140),
    .X(_0170_));
 sky130_fd_sc_hd__and2_1 _1562_ (.A(net406),
    .B(net140),
    .X(_0171_));
 sky130_fd_sc_hd__and2_1 _1563_ (.A(net407),
    .B(net140),
    .X(_0172_));
 sky130_fd_sc_hd__nor2_4 _1564_ (.A(net313),
    .B(_0493_),
    .Y(_0505_));
 sky130_fd_sc_hd__clkbuf_4 _1565_ (.A(net314),
    .X(_0506_));
 sky130_fd_sc_hd__nor2_4 _1566_ (.A(_0521_),
    .B(net314),
    .Y(_0507_));
 sky130_fd_sc_hd__clkbuf_4 _1567_ (.A(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__a22o_1 _1568_ (.A1(net300),
    .A2(_0506_),
    .B1(_0508_),
    .B2(net33),
    .X(_0173_));
 sky130_fd_sc_hd__a22o_1 _1569_ (.A1(net294),
    .A2(_0506_),
    .B1(_0508_),
    .B2(net44),
    .X(_0174_));
 sky130_fd_sc_hd__a22o_1 _1570_ (.A1(net290),
    .A2(_0506_),
    .B1(_0508_),
    .B2(net55),
    .X(_0175_));
 sky130_fd_sc_hd__a22o_1 _1571_ (.A1(net292),
    .A2(_0506_),
    .B1(_0508_),
    .B2(net58),
    .X(_0176_));
 sky130_fd_sc_hd__a22o_1 _1572_ (.A1(\register_file.write_data[4] ),
    .A2(_0506_),
    .B1(_0508_),
    .B2(net389),
    .X(_0177_));
 sky130_fd_sc_hd__a22o_1 _1573_ (.A1(\register_file.write_data[5] ),
    .A2(_0506_),
    .B1(_0508_),
    .B2(net488),
    .X(_0178_));
 sky130_fd_sc_hd__a22o_1 _1574_ (.A1(net482),
    .A2(_0506_),
    .B1(_0508_),
    .B2(net366),
    .X(_0179_));
 sky130_fd_sc_hd__a22o_1 _1575_ (.A1(net481),
    .A2(_0506_),
    .B1(_0508_),
    .B2(net368),
    .X(_0180_));
 sky130_fd_sc_hd__a22o_1 _1576_ (.A1(net296),
    .A2(_0506_),
    .B1(_0508_),
    .B2(net63),
    .X(_0181_));
 sky130_fd_sc_hd__a22o_1 _1577_ (.A1(net302),
    .A2(_0506_),
    .B1(_0508_),
    .B2(net64),
    .X(_0182_));
 sky130_fd_sc_hd__a22o_1 _1578_ (.A1(net210),
    .A2(_0506_),
    .B1(_0508_),
    .B2(net270),
    .X(_0183_));
 sky130_fd_sc_hd__a22o_1 _1579_ (.A1(net218),
    .A2(_0506_),
    .B1(_0508_),
    .B2(net276),
    .X(_0184_));
 sky130_fd_sc_hd__clkbuf_4 _1580_ (.A(net314),
    .X(_0509_));
 sky130_fd_sc_hd__clkbuf_4 _1581_ (.A(_0507_),
    .X(_0510_));
 sky130_fd_sc_hd__a22o_1 _1582_ (.A1(net212),
    .A2(_0509_),
    .B1(_0510_),
    .B2(net272),
    .X(_0185_));
 sky130_fd_sc_hd__a22o_1 _1583_ (.A1(net220),
    .A2(_0509_),
    .B1(_0510_),
    .B2(net274),
    .X(_0186_));
 sky130_fd_sc_hd__a22o_1 _1584_ (.A1(net208),
    .A2(_0509_),
    .B1(_0510_),
    .B2(net262),
    .X(_0187_));
 sky130_fd_sc_hd__a22o_1 _1585_ (.A1(net204),
    .A2(_0509_),
    .B1(_0510_),
    .B2(net256),
    .X(_0188_));
 sky130_fd_sc_hd__a22o_1 _1586_ (.A1(net206),
    .A2(_0509_),
    .B1(_0510_),
    .B2(net254),
    .X(_0189_));
 sky130_fd_sc_hd__a22o_1 _1587_ (.A1(net214),
    .A2(_0509_),
    .B1(_0510_),
    .B2(net268),
    .X(_0190_));
 sky130_fd_sc_hd__a22o_1 _1588_ (.A1(net216),
    .A2(_0509_),
    .B1(_0510_),
    .B2(net266),
    .X(_0191_));
 sky130_fd_sc_hd__a22o_1 _1589_ (.A1(net202),
    .A2(_0509_),
    .B1(_0510_),
    .B2(net252),
    .X(_0192_));
 sky130_fd_sc_hd__a22o_1 _1590_ (.A1(net228),
    .A2(_0509_),
    .B1(_0510_),
    .B2(net320),
    .X(_0193_));
 sky130_fd_sc_hd__a22o_1 _1591_ (.A1(net226),
    .A2(_0509_),
    .B1(_0510_),
    .B2(net316),
    .X(_0194_));
 sky130_fd_sc_hd__a22o_1 _1592_ (.A1(net224),
    .A2(_0509_),
    .B1(_0510_),
    .B2(net304),
    .X(_0195_));
 sky130_fd_sc_hd__a22o_1 _1593_ (.A1(net222),
    .A2(_0509_),
    .B1(_0510_),
    .B2(net306),
    .X(_0196_));
 sky130_fd_sc_hd__a22o_1 _1594_ (.A1(net282),
    .A2(net314),
    .B1(_0507_),
    .B2(net318),
    .X(_0197_));
 sky130_fd_sc_hd__a22o_1 _1595_ (.A1(net278),
    .A2(net314),
    .B1(_0507_),
    .B2(net50),
    .X(_0198_));
 sky130_fd_sc_hd__a22o_1 _1596_ (.A1(net280),
    .A2(net314),
    .B1(_0507_),
    .B2(net349),
    .X(_0199_));
 sky130_fd_sc_hd__a22o_1 _1597_ (.A1(net494),
    .A2(net314),
    .B1(_0507_),
    .B2(net347),
    .X(_0200_));
 sky130_fd_sc_hd__a22o_1 _1598_ (.A1(net351),
    .A2(net314),
    .B1(_0507_),
    .B2(net357),
    .X(_0201_));
 sky130_fd_sc_hd__a22o_1 _1599_ (.A1(net341),
    .A2(net314),
    .B1(_0507_),
    .B2(net343),
    .X(_0202_));
 sky130_fd_sc_hd__a22o_1 _1600_ (.A1(net372),
    .A2(net314),
    .B1(_0507_),
    .B2(net56),
    .X(_0203_));
 sky130_fd_sc_hd__a22o_1 _1601_ (.A1(net378),
    .A2(net314),
    .B1(_0507_),
    .B2(net57),
    .X(_0204_));
 sky130_fd_sc_hd__nor2_4 _1602_ (.A(net308),
    .B(_0493_),
    .Y(_0511_));
 sky130_fd_sc_hd__clkbuf_4 _1603_ (.A(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__nor2_4 _1604_ (.A(_0521_),
    .B(net309),
    .Y(_0513_));
 sky130_fd_sc_hd__clkbuf_4 _1605_ (.A(_0513_),
    .X(_0514_));
 sky130_fd_sc_hd__a22o_1 _1606_ (.A1(net300),
    .A2(_0512_),
    .B1(_0514_),
    .B2(net483),
    .X(_0205_));
 sky130_fd_sc_hd__a22o_1 _1607_ (.A1(net294),
    .A2(_0512_),
    .B1(_0514_),
    .B2(net478),
    .X(_0206_));
 sky130_fd_sc_hd__a22o_1 _1608_ (.A1(net290),
    .A2(_0512_),
    .B1(_0514_),
    .B2(net501),
    .X(_0207_));
 sky130_fd_sc_hd__a22o_1 _1609_ (.A1(net292),
    .A2(_0512_),
    .B1(_0514_),
    .B2(net486),
    .X(_0208_));
 sky130_fd_sc_hd__a22o_1 _1610_ (.A1(\register_file.write_data[4] ),
    .A2(_0512_),
    .B1(_0514_),
    .B2(net477),
    .X(_0209_));
 sky130_fd_sc_hd__a22o_1 _1611_ (.A1(\register_file.write_data[5] ),
    .A2(_0512_),
    .B1(_0514_),
    .B2(net264),
    .X(_0210_));
 sky130_fd_sc_hd__a22o_1 _1612_ (.A1(\register_file.write_data[6] ),
    .A2(_0512_),
    .B1(_0514_),
    .B2(net260),
    .X(_0211_));
 sky130_fd_sc_hd__a22o_1 _1613_ (.A1(\register_file.write_data[7] ),
    .A2(_0512_),
    .B1(_0514_),
    .B2(net258),
    .X(_0212_));
 sky130_fd_sc_hd__a22o_1 _1614_ (.A1(net296),
    .A2(_0512_),
    .B1(_0514_),
    .B2(net284),
    .X(_0213_));
 sky130_fd_sc_hd__a22o_1 _1615_ (.A1(net302),
    .A2(_0512_),
    .B1(_0514_),
    .B2(net298),
    .X(_0214_));
 sky130_fd_sc_hd__a22o_1 _1616_ (.A1(net210),
    .A2(_0512_),
    .B1(_0514_),
    .B2(net2),
    .X(_0215_));
 sky130_fd_sc_hd__a22o_1 _1617_ (.A1(net218),
    .A2(_0512_),
    .B1(_0514_),
    .B2(net3),
    .X(_0216_));
 sky130_fd_sc_hd__clkbuf_4 _1618_ (.A(_0511_),
    .X(_0515_));
 sky130_fd_sc_hd__clkbuf_4 _1619_ (.A(_0513_),
    .X(_0516_));
 sky130_fd_sc_hd__a22o_1 _1620_ (.A1(net212),
    .A2(_0515_),
    .B1(_0516_),
    .B2(net4),
    .X(_0217_));
 sky130_fd_sc_hd__a22o_1 _1621_ (.A1(net220),
    .A2(_0515_),
    .B1(_0516_),
    .B2(net5),
    .X(_0218_));
 sky130_fd_sc_hd__a22o_1 _1622_ (.A1(net208),
    .A2(_0515_),
    .B1(_0516_),
    .B2(net6),
    .X(_0219_));
 sky130_fd_sc_hd__a22o_1 _1623_ (.A1(net204),
    .A2(_0515_),
    .B1(_0516_),
    .B2(net7),
    .X(_0220_));
 sky130_fd_sc_hd__a22o_1 _1624_ (.A1(net206),
    .A2(_0515_),
    .B1(_0516_),
    .B2(net8),
    .X(_0221_));
 sky130_fd_sc_hd__a22o_1 _1625_ (.A1(net214),
    .A2(_0515_),
    .B1(_0516_),
    .B2(net9),
    .X(_0222_));
 sky130_fd_sc_hd__a22o_1 _1626_ (.A1(net216),
    .A2(_0515_),
    .B1(_0516_),
    .B2(net10),
    .X(_0223_));
 sky130_fd_sc_hd__a22o_1 _1627_ (.A1(net202),
    .A2(_0515_),
    .B1(_0516_),
    .B2(net11),
    .X(_0224_));
 sky130_fd_sc_hd__a22o_1 _1628_ (.A1(net228),
    .A2(_0515_),
    .B1(_0516_),
    .B2(net13),
    .X(_0225_));
 sky130_fd_sc_hd__a22o_1 _1629_ (.A1(net226),
    .A2(_0515_),
    .B1(_0516_),
    .B2(net14),
    .X(_0226_));
 sky130_fd_sc_hd__a22o_1 _1630_ (.A1(net224),
    .A2(_0515_),
    .B1(_0516_),
    .B2(net15),
    .X(_0227_));
 sky130_fd_sc_hd__a22o_1 _1631_ (.A1(net222),
    .A2(_0515_),
    .B1(_0516_),
    .B2(net16),
    .X(_0228_));
 sky130_fd_sc_hd__a22o_1 _1632_ (.A1(net282),
    .A2(net309),
    .B1(_0513_),
    .B2(net17),
    .X(_0229_));
 sky130_fd_sc_hd__a22o_1 _1633_ (.A1(net278),
    .A2(net309),
    .B1(_0513_),
    .B2(net311),
    .X(_0230_));
 sky130_fd_sc_hd__a22o_1 _1634_ (.A1(net280),
    .A2(net309),
    .B1(_0513_),
    .B2(net409),
    .X(_0231_));
 sky130_fd_sc_hd__a22o_1 _1635_ (.A1(net494),
    .A2(net309),
    .B1(_0513_),
    .B2(net339),
    .X(_0232_));
 sky130_fd_sc_hd__a22o_1 _1636_ (.A1(net351),
    .A2(net309),
    .B1(_0513_),
    .B2(net355),
    .X(_0233_));
 sky130_fd_sc_hd__a22o_1 _1637_ (.A1(net341),
    .A2(net309),
    .B1(_0513_),
    .B2(net345),
    .X(_0234_));
 sky130_fd_sc_hd__a22o_1 _1638_ (.A1(net372),
    .A2(net309),
    .B1(_0513_),
    .B2(net353),
    .X(_0235_));
 sky130_fd_sc_hd__a22o_1 _1639_ (.A1(net378),
    .A2(net309),
    .B1(_0513_),
    .B2(net487),
    .X(_0236_));
 sky130_fd_sc_hd__and2_1 _1640_ (.A(_0442_),
    .B(net510),
    .X(_0237_));
 sky130_fd_sc_hd__inv_2 _1641_ (.A(_0522_),
    .Y(_0238_));
 sky130_fd_sc_hd__nor2_1 _1642_ (.A(net337),
    .B(_0521_),
    .Y(_0239_));
 sky130_fd_sc_hd__and3_1 _1643_ (.A(_0441_),
    .B(_0411_),
    .C(net483),
    .X(_0240_));
 sky130_fd_sc_hd__and3_1 _1644_ (.A(_0441_),
    .B(_0411_),
    .C(net478),
    .X(_0241_));
 sky130_fd_sc_hd__and3_1 _1645_ (.A(_0441_),
    .B(_0411_),
    .C(net501),
    .X(_0242_));
 sky130_fd_sc_hd__and3_1 _1646_ (.A(_0441_),
    .B(_0411_),
    .C(net486),
    .X(_0243_));
 sky130_fd_sc_hd__and3_1 _1647_ (.A(_0441_),
    .B(_0411_),
    .C(net477),
    .X(_0244_));
 sky130_fd_sc_hd__and3_1 _1648_ (.A(_0441_),
    .B(_0411_),
    .C(net264),
    .X(_0245_));
 sky130_fd_sc_hd__and3_1 _1649_ (.A(_0441_),
    .B(_0411_),
    .C(net260),
    .X(_0246_));
 sky130_fd_sc_hd__and3_1 _1650_ (.A(_0441_),
    .B(_0411_),
    .C(net258),
    .X(_0247_));
 sky130_fd_sc_hd__and3_1 _1651_ (.A(_0441_),
    .B(_0411_),
    .C(net284),
    .X(_0248_));
 sky130_fd_sc_hd__and3_1 _1652_ (.A(_0441_),
    .B(_0411_),
    .C(net298),
    .X(_0249_));
 sky130_fd_sc_hd__and3_1 _1653_ (.A(_0441_),
    .B(_0411_),
    .C(net361),
    .X(_0250_));
 sky130_fd_sc_hd__clkbuf_2 _1654_ (.A(net337),
    .X(_0517_));
 sky130_fd_sc_hd__buf_1 _1655_ (.A(_0519_),
    .X(_0518_));
 sky130_fd_sc_hd__and3_1 _1656_ (.A(_0517_),
    .B(_0518_),
    .C(net362),
    .X(_0251_));
 sky130_fd_sc_hd__and3_1 _1657_ (.A(_0517_),
    .B(_0518_),
    .C(net365),
    .X(_0252_));
 sky130_fd_sc_hd__and3_1 _1658_ (.A(_0517_),
    .B(_0518_),
    .C(net5),
    .X(_0253_));
 sky130_fd_sc_hd__and3_1 _1659_ (.A(_0517_),
    .B(_0518_),
    .C(net6),
    .X(_0254_));
 sky130_fd_sc_hd__and3_1 _1660_ (.A(_0517_),
    .B(_0518_),
    .C(net7),
    .X(_0255_));
 sky130_fd_sc_hd__and3_1 _1661_ (.A(_0517_),
    .B(_0518_),
    .C(net8),
    .X(_0256_));
 sky130_fd_sc_hd__and3_1 _1662_ (.A(_0517_),
    .B(_0518_),
    .C(net363),
    .X(_0257_));
 sky130_fd_sc_hd__and3_1 _1663_ (.A(_0517_),
    .B(_0518_),
    .C(net10),
    .X(_0258_));
 sky130_fd_sc_hd__and3_1 _1664_ (.A(_0517_),
    .B(_0518_),
    .C(net519),
    .X(_0259_));
 sky130_fd_sc_hd__and3_1 _1665_ (.A(_0517_),
    .B(_0518_),
    .C(net364),
    .X(_0260_));
 sky130_fd_sc_hd__and3_1 _1666_ (.A(_0517_),
    .B(_0518_),
    .C(net14),
    .X(_0261_));
 sky130_fd_sc_hd__and3_1 _1667_ (.A(_0517_),
    .B(_0518_),
    .C(net524),
    .X(_0262_));
 sky130_fd_sc_hd__and3_1 _1668_ (.A(net337),
    .B(_0592_),
    .C(net16),
    .X(_0263_));
 sky130_fd_sc_hd__and3_1 _1669_ (.A(net337),
    .B(_0592_),
    .C(net535),
    .X(_0264_));
 sky130_fd_sc_hd__and3_1 _1670_ (.A(net337),
    .B(_0592_),
    .C(net311),
    .X(_0265_));
 sky130_fd_sc_hd__and3_1 _1671_ (.A(net337),
    .B(_0592_),
    .C(net409),
    .X(_0266_));
 sky130_fd_sc_hd__and3_1 _1672_ (.A(net337),
    .B(_0592_),
    .C(net339),
    .X(_0267_));
 sky130_fd_sc_hd__and3_1 _1673_ (.A(net337),
    .B(_0592_),
    .C(net355),
    .X(_0268_));
 sky130_fd_sc_hd__and3_1 _1674_ (.A(net337),
    .B(_0592_),
    .C(net345),
    .X(_0269_));
 sky130_fd_sc_hd__and3_1 _1675_ (.A(net337),
    .B(_0592_),
    .C(net353),
    .X(_0270_));
 sky130_fd_sc_hd__and3_1 _1676_ (.A(net337),
    .B(_0592_),
    .C(net487),
    .X(_0271_));
 sky130_fd_sc_hd__and2_1 _1677_ (.A(net490),
    .B(_0239_),
    .X(_0272_));
 sky130_fd_sc_hd__and2_1 _1678_ (.A(net408),
    .B(_0239_),
    .X(_0273_));
 sky130_fd_sc_hd__and2_1 _1679_ (.A(net404),
    .B(_0239_),
    .X(_0274_));
 sky130_fd_sc_hd__nor2_1 _1680_ (.A(net434),
    .B(net473),
    .Y(_0275_));
 sky130_fd_sc_hd__nor2b_1 _1681_ (.A(_0443_),
    .B_N(_0275_),
    .Y(_0276_));
 sky130_fd_sc_hd__nor2b_1 _1682_ (.A(net330),
    .B_N(_0275_),
    .Y(_0277_));
 sky130_fd_sc_hd__nor2_1 _1683_ (.A(_0440_),
    .B(_0443_),
    .Y(_0278_));
 sky130_fd_sc_hd__dfxtp_2 _1684_ (.CLK(clknet_leaf_20_clk),
    .D(_0001_),
    .Q(\register_file.write_data[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1685_ (.CLK(clknet_leaf_20_clk),
    .D(_0002_),
    .Q(\register_file.write_data[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1686_ (.CLK(clknet_leaf_20_clk),
    .D(_0003_),
    .Q(\register_file.write_data[2] ));
 sky130_fd_sc_hd__dfxtp_2 _1687_ (.CLK(clknet_leaf_20_clk),
    .D(_0004_),
    .Q(\register_file.write_data[3] ));
 sky130_fd_sc_hd__dfxtp_2 _1688_ (.CLK(clknet_leaf_0_clk),
    .D(net231),
    .Q(\register_file.write_data[4] ));
 sky130_fd_sc_hd__dfxtp_2 _1689_ (.CLK(clknet_leaf_0_clk),
    .D(_0006_),
    .Q(\register_file.write_data[5] ));
 sky130_fd_sc_hd__dfxtp_2 _1690_ (.CLK(clknet_leaf_0_clk),
    .D(net197),
    .Q(\register_file.write_data[6] ));
 sky130_fd_sc_hd__dfxtp_2 _1691_ (.CLK(clknet_leaf_0_clk),
    .D(net199),
    .Q(\register_file.write_data[7] ));
 sky130_fd_sc_hd__dfxtp_2 _1692_ (.CLK(clknet_leaf_19_clk),
    .D(_0009_),
    .Q(\register_file.write_data[8] ));
 sky130_fd_sc_hd__dfxtp_2 _1693_ (.CLK(clknet_leaf_19_clk),
    .D(_0010_),
    .Q(\register_file.write_data[9] ));
 sky130_fd_sc_hd__dfxtp_2 _1694_ (.CLK(clknet_leaf_17_clk),
    .D(_0011_),
    .Q(\register_file.write_data[10] ));
 sky130_fd_sc_hd__dfxtp_2 _1695_ (.CLK(clknet_leaf_3_clk),
    .D(_0012_),
    .Q(\register_file.write_data[11] ));
 sky130_fd_sc_hd__dfxtp_2 _1696_ (.CLK(clknet_leaf_3_clk),
    .D(_0013_),
    .Q(\register_file.write_data[12] ));
 sky130_fd_sc_hd__dfxtp_2 _1697_ (.CLK(clknet_leaf_3_clk),
    .D(_0014_),
    .Q(\register_file.write_data[13] ));
 sky130_fd_sc_hd__dfxtp_2 _1698_ (.CLK(clknet_leaf_3_clk),
    .D(_0015_),
    .Q(\register_file.write_data[14] ));
 sky130_fd_sc_hd__dfxtp_2 _1699_ (.CLK(clknet_leaf_3_clk),
    .D(_0016_),
    .Q(\register_file.write_data[15] ));
 sky130_fd_sc_hd__dfxtp_2 _1700_ (.CLK(clknet_leaf_3_clk),
    .D(net377),
    .Q(\register_file.write_data[16] ));
 sky130_fd_sc_hd__dfxtp_2 _1701_ (.CLK(clknet_leaf_3_clk),
    .D(net375),
    .Q(\register_file.write_data[17] ));
 sky130_fd_sc_hd__dfxtp_2 _1702_ (.CLK(clknet_leaf_3_clk),
    .D(net381),
    .Q(\register_file.write_data[18] ));
 sky130_fd_sc_hd__dfxtp_2 _1703_ (.CLK(clknet_leaf_3_clk),
    .D(net371),
    .Q(\register_file.write_data[19] ));
 sky130_fd_sc_hd__dfxtp_2 _1704_ (.CLK(clknet_leaf_5_clk),
    .D(net336),
    .Q(\register_file.write_data[20] ));
 sky130_fd_sc_hd__dfxtp_2 _1705_ (.CLK(clknet_leaf_5_clk),
    .D(net323),
    .Q(\register_file.write_data[21] ));
 sky130_fd_sc_hd__dfxtp_2 _1706_ (.CLK(clknet_leaf_5_clk),
    .D(net327),
    .Q(\register_file.write_data[22] ));
 sky130_fd_sc_hd__dfxtp_2 _1707_ (.CLK(clknet_leaf_5_clk),
    .D(net329),
    .Q(\register_file.write_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 _1708_ (.CLK(clknet_leaf_5_clk),
    .D(_0025_),
    .Q(\register_file.write_data[24] ));
 sky130_fd_sc_hd__dfxtp_1 _1709_ (.CLK(clknet_leaf_5_clk),
    .D(_0026_),
    .Q(\register_file.write_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 _1710_ (.CLK(clknet_leaf_5_clk),
    .D(net325),
    .Q(\register_file.write_data[26] ));
 sky130_fd_sc_hd__dfxtp_1 _1711_ (.CLK(clknet_leaf_8_clk),
    .D(net201),
    .Q(\register_file.write_data[27] ));
 sky130_fd_sc_hd__dfxtp_2 _1712_ (.CLK(clknet_leaf_10_clk),
    .D(_0029_),
    .Q(\register_file.write_data[28] ));
 sky130_fd_sc_hd__dfxtp_2 _1713_ (.CLK(clknet_leaf_10_clk),
    .D(_0030_),
    .Q(\register_file.write_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 _1714_ (.CLK(clknet_leaf_10_clk),
    .D(_0031_),
    .Q(\register_file.write_data[30] ));
 sky130_fd_sc_hd__dfxtp_1 _1715_ (.CLK(clknet_leaf_10_clk),
    .D(_0032_),
    .Q(\register_file.write_data[31] ));
 sky130_fd_sc_hd__dfxtp_1 _1716_ (.CLK(clknet_leaf_20_clk),
    .D(net509),
    .Q(\ex_mem_alu_result[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1717_ (.CLK(clknet_leaf_20_clk),
    .D(net529),
    .Q(\ex_mem_alu_result[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1718_ (.CLK(clknet_leaf_20_clk),
    .D(net532),
    .Q(\dmem.address[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1719_ (.CLK(clknet_leaf_20_clk),
    .D(net523),
    .Q(\dmem.address[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1720_ (.CLK(clknet_leaf_20_clk),
    .D(_0037_),
    .Q(\dmem.address[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1721_ (.CLK(clknet_leaf_0_clk),
    .D(net400),
    .Q(\dmem.address[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1722_ (.CLK(clknet_leaf_19_clk),
    .D(_0039_),
    .Q(\dmem.address[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1723_ (.CLK(clknet_leaf_19_clk),
    .D(_0040_),
    .Q(\dmem.address[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1724_ (.CLK(clknet_leaf_17_clk),
    .D(_0041_),
    .Q(\dmem.address[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1725_ (.CLK(clknet_leaf_17_clk),
    .D(_0042_),
    .Q(\dmem.address[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1726_ (.CLK(clknet_leaf_17_clk),
    .D(_0043_),
    .Q(\dmem.address[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1727_ (.CLK(clknet_leaf_17_clk),
    .D(_0044_),
    .Q(\dmem.address[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1728_ (.CLK(clknet_leaf_17_clk),
    .D(_0045_),
    .Q(\dmem.address[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1729_ (.CLK(clknet_leaf_17_clk),
    .D(_0046_),
    .Q(\dmem.address[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1730_ (.CLK(clknet_leaf_4_clk),
    .D(_0047_),
    .Q(\dmem.address[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1731_ (.CLK(clknet_leaf_4_clk),
    .D(_0048_),
    .Q(\dmem.address[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1732_ (.CLK(clknet_leaf_4_clk),
    .D(_0049_),
    .Q(\dmem.address[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1733_ (.CLK(clknet_leaf_4_clk),
    .D(_0050_),
    .Q(\dmem.address[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1734_ (.CLK(clknet_leaf_4_clk),
    .D(_0051_),
    .Q(\dmem.address[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1735_ (.CLK(clknet_leaf_4_clk),
    .D(_0052_),
    .Q(\dmem.address[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1736_ (.CLK(clknet_leaf_4_clk),
    .D(_0053_),
    .Q(\dmem.address[20] ));
 sky130_fd_sc_hd__dfxtp_1 _1737_ (.CLK(clknet_leaf_4_clk),
    .D(_0054_),
    .Q(\dmem.address[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1738_ (.CLK(clknet_leaf_4_clk),
    .D(_0055_),
    .Q(\dmem.address[22] ));
 sky130_fd_sc_hd__dfxtp_1 _1739_ (.CLK(clknet_leaf_4_clk),
    .D(_0056_),
    .Q(\dmem.address[23] ));
 sky130_fd_sc_hd__dfxtp_1 _1740_ (.CLK(clknet_leaf_5_clk),
    .D(_0057_),
    .Q(\dmem.address[24] ));
 sky130_fd_sc_hd__dfxtp_1 _1741_ (.CLK(clknet_leaf_5_clk),
    .D(_0058_),
    .Q(\dmem.address[25] ));
 sky130_fd_sc_hd__dfxtp_1 _1742_ (.CLK(clknet_leaf_11_clk),
    .D(_0059_),
    .Q(\dmem.address[26] ));
 sky130_fd_sc_hd__dfxtp_1 _1743_ (.CLK(clknet_leaf_11_clk),
    .D(_0060_),
    .Q(\dmem.address[27] ));
 sky130_fd_sc_hd__dfxtp_1 _1744_ (.CLK(clknet_leaf_10_clk),
    .D(net496),
    .Q(\dmem.address[28] ));
 sky130_fd_sc_hd__dfxtp_1 _1745_ (.CLK(clknet_leaf_10_clk),
    .D(_0062_),
    .Q(\dmem.address[29] ));
 sky130_fd_sc_hd__dfxtp_1 _1746_ (.CLK(clknet_leaf_10_clk),
    .D(_0063_),
    .Q(\dmem.address[30] ));
 sky130_fd_sc_hd__dfxtp_1 _1747_ (.CLK(clknet_leaf_10_clk),
    .D(_0064_),
    .Q(\dmem.address[31] ));
 sky130_fd_sc_hd__dfxtp_2 _1748_ (.CLK(clknet_leaf_9_clk),
    .D(_0065_),
    .Q(mem_wb_valid));
 sky130_fd_sc_hd__dfxtp_1 _1749_ (.CLK(clknet_leaf_9_clk),
    .D(_0066_),
    .Q(ex_mem_valid));
 sky130_fd_sc_hd__dfxtp_2 _1750_ (.CLK(clknet_leaf_19_clk),
    .D(_0067_),
    .Q(\forwarding_unit.rd_wb[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1751_ (.CLK(clknet_leaf_19_clk),
    .D(_0068_),
    .Q(\forwarding_unit.rd_wb[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1752_ (.CLK(clknet_leaf_16_clk),
    .D(_0069_),
    .Q(net101));
 sky130_fd_sc_hd__dfxtp_1 _1753_ (.CLK(clknet_leaf_20_clk),
    .D(_0070_),
    .Q(\forwarding_unit.rs1_ex[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1754_ (.CLK(clknet_leaf_19_clk),
    .D(_0071_),
    .Q(\forwarding_unit.rs2_ex[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1755_ (.CLK(clknet_leaf_19_clk),
    .D(_0072_),
    .Q(\forwarding_unit.rs2_ex[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1756_ (.CLK(clknet_leaf_19_clk),
    .D(_0073_),
    .Q(\forwarding_unit.rs2_ex[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1757_ (.CLK(clknet_leaf_19_clk),
    .D(_0074_),
    .Q(\id_ex_rd_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1758_ (.CLK(clknet_leaf_9_clk),
    .D(_0075_),
    .Q(id_ex_valid));
 sky130_fd_sc_hd__dfxtp_1 _1759_ (.CLK(clknet_leaf_9_clk),
    .D(_0000_),
    .Q(if_id_valid));
 sky130_fd_sc_hd__dfxtp_1 _1760_ (.CLK(clknet_leaf_18_clk),
    .D(net334),
    .Q(\forwarding_unit.rd_mem[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1761_ (.CLK(clknet_leaf_19_clk),
    .D(_0077_),
    .Q(\forwarding_unit.rd_mem[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1762_ (.CLK(clknet_leaf_19_clk),
    .D(_0078_),
    .Q(\forwarding_unit.reg_write_wb ));
 sky130_fd_sc_hd__dfxtp_4 _1763_ (.CLK(clknet_leaf_15_clk),
    .D(_0079_),
    .Q(net125));
 sky130_fd_sc_hd__dfxtp_2 _1764_ (.CLK(clknet_leaf_16_clk),
    .D(_0080_),
    .Q(net128));
 sky130_fd_sc_hd__dfxtp_2 _1765_ (.CLK(clknet_leaf_15_clk),
    .D(net332),
    .Q(net129));
 sky130_fd_sc_hd__dfxtp_1 _1766_ (.CLK(clknet_leaf_15_clk),
    .D(net403),
    .Q(net130));
 sky130_fd_sc_hd__dfxtp_1 _1767_ (.CLK(clknet_leaf_14_clk),
    .D(_0083_),
    .Q(net131));
 sky130_fd_sc_hd__dfxtp_1 _1768_ (.CLK(clknet_leaf_14_clk),
    .D(_0084_),
    .Q(net132));
 sky130_fd_sc_hd__dfxtp_1 _1769_ (.CLK(clknet_leaf_14_clk),
    .D(net493),
    .Q(net133));
 sky130_fd_sc_hd__dfxtp_1 _1770_ (.CLK(clknet_leaf_14_clk),
    .D(_0086_),
    .Q(net134));
 sky130_fd_sc_hd__dfxtp_1 _1771_ (.CLK(clknet_leaf_14_clk),
    .D(net504),
    .Q(net105));
 sky130_fd_sc_hd__dfxtp_1 _1772_ (.CLK(clknet_leaf_14_clk),
    .D(_0088_),
    .Q(net106));
 sky130_fd_sc_hd__dfxtp_1 _1773_ (.CLK(clknet_leaf_14_clk),
    .D(_0089_),
    .Q(net107));
 sky130_fd_sc_hd__dfxtp_1 _1774_ (.CLK(clknet_leaf_14_clk),
    .D(_0090_),
    .Q(net108));
 sky130_fd_sc_hd__dfxtp_1 _1775_ (.CLK(clknet_leaf_13_clk),
    .D(net417),
    .Q(net109));
 sky130_fd_sc_hd__dfxtp_1 _1776_ (.CLK(clknet_leaf_13_clk),
    .D(net515),
    .Q(net110));
 sky130_fd_sc_hd__dfxtp_1 _1777_ (.CLK(clknet_leaf_13_clk),
    .D(net468),
    .Q(net111));
 sky130_fd_sc_hd__dfxtp_1 _1778_ (.CLK(clknet_leaf_13_clk),
    .D(net452),
    .Q(net112));
 sky130_fd_sc_hd__dfxtp_1 _1779_ (.CLK(clknet_leaf_13_clk),
    .D(_0095_),
    .Q(net113));
 sky130_fd_sc_hd__dfxtp_1 _1780_ (.CLK(clknet_leaf_13_clk),
    .D(net465),
    .Q(net114));
 sky130_fd_sc_hd__dfxtp_1 _1781_ (.CLK(clknet_leaf_13_clk),
    .D(net448),
    .Q(net115));
 sky130_fd_sc_hd__dfxtp_1 _1782_ (.CLK(clknet_leaf_13_clk),
    .D(_0098_),
    .Q(net116));
 sky130_fd_sc_hd__dfxtp_1 _1783_ (.CLK(clknet_leaf_12_clk),
    .D(net428),
    .Q(net117));
 sky130_fd_sc_hd__dfxtp_1 _1784_ (.CLK(clknet_leaf_12_clk),
    .D(net450),
    .Q(net118));
 sky130_fd_sc_hd__dfxtp_1 _1785_ (.CLK(clknet_leaf_12_clk),
    .D(net513),
    .Q(net119));
 sky130_fd_sc_hd__dfxtp_1 _1786_ (.CLK(clknet_leaf_12_clk),
    .D(net462),
    .Q(net120));
 sky130_fd_sc_hd__dfxtp_1 _1787_ (.CLK(clknet_leaf_12_clk),
    .D(net456),
    .Q(net121));
 sky130_fd_sc_hd__dfxtp_1 _1788_ (.CLK(clknet_leaf_12_clk),
    .D(_0104_),
    .Q(net122));
 sky130_fd_sc_hd__dfxtp_1 _1789_ (.CLK(clknet_leaf_12_clk),
    .D(net476),
    .Q(net123));
 sky130_fd_sc_hd__dfxtp_1 _1790_ (.CLK(clknet_leaf_12_clk),
    .D(net485),
    .Q(net124));
 sky130_fd_sc_hd__dfxtp_1 _1791_ (.CLK(clknet_leaf_12_clk),
    .D(net480),
    .Q(net126));
 sky130_fd_sc_hd__dfxtp_1 _1792_ (.CLK(clknet_leaf_12_clk),
    .D(_0108_),
    .Q(net127));
 sky130_fd_sc_hd__dfxtp_1 _1793_ (.CLK(clknet_leaf_7_clk),
    .D(_0109_),
    .Q(net65));
 sky130_fd_sc_hd__dfxtp_1 _1794_ (.CLK(clknet_leaf_7_clk),
    .D(_0110_),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_1 _1795_ (.CLK(clknet_leaf_7_clk),
    .D(_0111_),
    .Q(net87));
 sky130_fd_sc_hd__dfxtp_1 _1796_ (.CLK(clknet_leaf_7_clk),
    .D(_0112_),
    .Q(net90));
 sky130_fd_sc_hd__dfxtp_1 _1797_ (.CLK(clknet_leaf_7_clk),
    .D(_0113_),
    .Q(net91));
 sky130_fd_sc_hd__dfxtp_1 _1798_ (.CLK(clknet_leaf_7_clk),
    .D(_0114_),
    .Q(net92));
 sky130_fd_sc_hd__dfxtp_1 _1799_ (.CLK(clknet_leaf_7_clk),
    .D(_0115_),
    .Q(net93));
 sky130_fd_sc_hd__dfxtp_1 _1800_ (.CLK(clknet_leaf_7_clk),
    .D(_0116_),
    .Q(net94));
 sky130_fd_sc_hd__dfxtp_1 _1801_ (.CLK(clknet_leaf_7_clk),
    .D(_0117_),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_1 _1802_ (.CLK(clknet_leaf_7_clk),
    .D(_0118_),
    .Q(net96));
 sky130_fd_sc_hd__dfxtp_1 _1803_ (.CLK(clknet_leaf_7_clk),
    .D(_0119_),
    .Q(net66));
 sky130_fd_sc_hd__dfxtp_1 _1804_ (.CLK(clknet_leaf_7_clk),
    .D(_0120_),
    .Q(net67));
 sky130_fd_sc_hd__dfxtp_1 _1805_ (.CLK(clknet_leaf_9_clk),
    .D(net241),
    .Q(net68));
 sky130_fd_sc_hd__dfxtp_1 _1806_ (.CLK(clknet_leaf_8_clk),
    .D(net247),
    .Q(net69));
 sky130_fd_sc_hd__dfxtp_1 _1807_ (.CLK(clknet_leaf_9_clk),
    .D(net235),
    .Q(net70));
 sky130_fd_sc_hd__dfxtp_1 _1808_ (.CLK(clknet_leaf_9_clk),
    .D(net239),
    .Q(net71));
 sky130_fd_sc_hd__dfxtp_1 _1809_ (.CLK(clknet_leaf_8_clk),
    .D(net237),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_1 _1810_ (.CLK(clknet_leaf_9_clk),
    .D(net243),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_1 _1811_ (.CLK(clknet_leaf_9_clk),
    .D(net245),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_1 _1812_ (.CLK(clknet_leaf_9_clk),
    .D(net233),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_1 _1813_ (.CLK(clknet_leaf_9_clk),
    .D(net289),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_1 _1814_ (.CLK(clknet_leaf_9_clk),
    .D(net287),
    .Q(net78));
 sky130_fd_sc_hd__dfxtp_1 _1815_ (.CLK(clknet_leaf_9_clk),
    .D(net249),
    .Q(net79));
 sky130_fd_sc_hd__dfxtp_1 _1816_ (.CLK(clknet_leaf_9_clk),
    .D(net251),
    .Q(net80));
 sky130_fd_sc_hd__dfxtp_1 _1817_ (.CLK(clknet_leaf_8_clk),
    .D(net283),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_1 _1818_ (.CLK(clknet_leaf_8_clk),
    .D(net279),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_1 _1819_ (.CLK(clknet_leaf_9_clk),
    .D(net281),
    .Q(net83));
 sky130_fd_sc_hd__dfxtp_1 _1820_ (.CLK(clknet_leaf_9_clk),
    .D(net470),
    .Q(net84));
 sky130_fd_sc_hd__dfxtp_1 _1821_ (.CLK(clknet_leaf_9_clk),
    .D(net352),
    .Q(net85));
 sky130_fd_sc_hd__dfxtp_1 _1822_ (.CLK(clknet_leaf_9_clk),
    .D(net342),
    .Q(net86));
 sky130_fd_sc_hd__dfxtp_1 _1823_ (.CLK(clknet_leaf_9_clk),
    .D(_0139_),
    .Q(net88));
 sky130_fd_sc_hd__dfxtp_1 _1824_ (.CLK(clknet_leaf_9_clk),
    .D(_0140_),
    .Q(net89));
 sky130_fd_sc_hd__dfxtp_1 _1825_ (.CLK(clknet_leaf_21_clk),
    .D(_0141_),
    .Q(\id_ex_rs2_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1826_ (.CLK(clknet_leaf_21_clk),
    .D(_0142_),
    .Q(\id_ex_rs2_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1827_ (.CLK(clknet_leaf_0_clk),
    .D(_0143_),
    .Q(\id_ex_rs2_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1828_ (.CLK(clknet_leaf_21_clk),
    .D(_0144_),
    .Q(\id_ex_rs2_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1829_ (.CLK(clknet_leaf_0_clk),
    .D(_0145_),
    .Q(\id_ex_rs2_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1830_ (.CLK(clknet_leaf_2_clk),
    .D(_0146_),
    .Q(\id_ex_rs2_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1831_ (.CLK(clknet_leaf_1_clk),
    .D(net367),
    .Q(\id_ex_rs2_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1832_ (.CLK(clknet_leaf_1_clk),
    .D(net369),
    .Q(\id_ex_rs2_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1833_ (.CLK(clknet_leaf_21_clk),
    .D(_0149_),
    .Q(\id_ex_rs2_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1834_ (.CLK(clknet_leaf_0_clk),
    .D(net384),
    .Q(\id_ex_rs2_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1835_ (.CLK(clknet_leaf_2_clk),
    .D(_0151_),
    .Q(\id_ex_rs2_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1836_ (.CLK(clknet_leaf_2_clk),
    .D(_0152_),
    .Q(\id_ex_rs2_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1837_ (.CLK(clknet_leaf_2_clk),
    .D(_0153_),
    .Q(\id_ex_rs2_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1838_ (.CLK(clknet_leaf_2_clk),
    .D(_0154_),
    .Q(\id_ex_rs2_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1839_ (.CLK(clknet_leaf_2_clk),
    .D(_0155_),
    .Q(\id_ex_rs2_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1840_ (.CLK(clknet_leaf_2_clk),
    .D(_0156_),
    .Q(\id_ex_rs2_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1841_ (.CLK(clknet_leaf_2_clk),
    .D(_0157_),
    .Q(\id_ex_rs2_data[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1842_ (.CLK(clknet_leaf_2_clk),
    .D(_0158_),
    .Q(\id_ex_rs2_data[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1843_ (.CLK(clknet_leaf_6_clk),
    .D(_0159_),
    .Q(\id_ex_rs2_data[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1844_ (.CLK(clknet_leaf_6_clk),
    .D(_0160_),
    .Q(\id_ex_rs2_data[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1845_ (.CLK(clknet_leaf_6_clk),
    .D(_0161_),
    .Q(\id_ex_rs2_data[20] ));
 sky130_fd_sc_hd__dfxtp_1 _1846_ (.CLK(clknet_leaf_6_clk),
    .D(_0162_),
    .Q(\id_ex_rs2_data[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1847_ (.CLK(clknet_leaf_6_clk),
    .D(_0163_),
    .Q(\id_ex_rs2_data[22] ));
 sky130_fd_sc_hd__dfxtp_1 _1848_ (.CLK(clknet_leaf_6_clk),
    .D(_0164_),
    .Q(\id_ex_rs2_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 _1849_ (.CLK(clknet_leaf_5_clk),
    .D(_0165_),
    .Q(\id_ex_rs2_data[24] ));
 sky130_fd_sc_hd__dfxtp_1 _1850_ (.CLK(clknet_leaf_5_clk),
    .D(_0166_),
    .Q(\id_ex_rs2_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 _1851_ (.CLK(clknet_leaf_8_clk),
    .D(net350),
    .Q(\id_ex_rs2_data[26] ));
 sky130_fd_sc_hd__dfxtp_1 _1852_ (.CLK(clknet_leaf_8_clk),
    .D(net348),
    .Q(\id_ex_rs2_data[27] ));
 sky130_fd_sc_hd__dfxtp_1 _1853_ (.CLK(clknet_leaf_8_clk),
    .D(_0169_),
    .Q(\id_ex_rs2_data[28] ));
 sky130_fd_sc_hd__dfxtp_1 _1854_ (.CLK(clknet_leaf_8_clk),
    .D(_0170_),
    .Q(\id_ex_rs2_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 _1855_ (.CLK(clknet_leaf_8_clk),
    .D(_0171_),
    .Q(\id_ex_rs2_data[30] ));
 sky130_fd_sc_hd__dfxtp_1 _1856_ (.CLK(clknet_leaf_8_clk),
    .D(_0172_),
    .Q(\id_ex_rs2_data[31] ));
 sky130_fd_sc_hd__dfxtp_2 _1857_ (.CLK(clknet_leaf_1_clk),
    .D(net301),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_2 _1858_ (.CLK(clknet_leaf_1_clk),
    .D(net295),
    .Q(net44));
 sky130_fd_sc_hd__dfxtp_2 _1859_ (.CLK(clknet_leaf_1_clk),
    .D(net291),
    .Q(net55));
 sky130_fd_sc_hd__dfxtp_2 _1860_ (.CLK(clknet_leaf_1_clk),
    .D(net293),
    .Q(net58));
 sky130_fd_sc_hd__dfxtp_2 _1861_ (.CLK(clknet_leaf_1_clk),
    .D(net390),
    .Q(net59));
 sky130_fd_sc_hd__dfxtp_1 _1862_ (.CLK(clknet_leaf_2_clk),
    .D(net489),
    .Q(net60));
 sky130_fd_sc_hd__dfxtp_1 _1863_ (.CLK(clknet_leaf_2_clk),
    .D(_0179_),
    .Q(net61));
 sky130_fd_sc_hd__dfxtp_1 _1864_ (.CLK(clknet_leaf_2_clk),
    .D(_0180_),
    .Q(net62));
 sky130_fd_sc_hd__dfxtp_1 _1865_ (.CLK(clknet_leaf_2_clk),
    .D(net297),
    .Q(net63));
 sky130_fd_sc_hd__dfxtp_1 _1866_ (.CLK(clknet_leaf_2_clk),
    .D(net303),
    .Q(net64));
 sky130_fd_sc_hd__dfxtp_1 _1867_ (.CLK(clknet_leaf_2_clk),
    .D(net271),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_1 _1868_ (.CLK(clknet_leaf_2_clk),
    .D(net277),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_1 _1869_ (.CLK(clknet_leaf_2_clk),
    .D(net273),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_1 _1870_ (.CLK(clknet_leaf_2_clk),
    .D(net275),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_1 _1871_ (.CLK(clknet_leaf_2_clk),
    .D(net263),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_1 _1872_ (.CLK(clknet_leaf_6_clk),
    .D(net257),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_1 _1873_ (.CLK(clknet_leaf_6_clk),
    .D(net255),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_1 _1874_ (.CLK(clknet_leaf_6_clk),
    .D(net269),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_1 _1875_ (.CLK(clknet_leaf_6_clk),
    .D(net267),
    .Q(net42));
 sky130_fd_sc_hd__dfxtp_1 _1876_ (.CLK(clknet_leaf_6_clk),
    .D(net253),
    .Q(net43));
 sky130_fd_sc_hd__dfxtp_1 _1877_ (.CLK(clknet_leaf_6_clk),
    .D(net321),
    .Q(net45));
 sky130_fd_sc_hd__dfxtp_1 _1878_ (.CLK(clknet_leaf_6_clk),
    .D(net317),
    .Q(net46));
 sky130_fd_sc_hd__dfxtp_1 _1879_ (.CLK(clknet_leaf_6_clk),
    .D(net305),
    .Q(net47));
 sky130_fd_sc_hd__dfxtp_1 _1880_ (.CLK(clknet_leaf_6_clk),
    .D(net307),
    .Q(net48));
 sky130_fd_sc_hd__dfxtp_1 _1881_ (.CLK(clknet_leaf_6_clk),
    .D(net319),
    .Q(net49));
 sky130_fd_sc_hd__dfxtp_1 _1882_ (.CLK(clknet_leaf_6_clk),
    .D(net315),
    .Q(net50));
 sky130_fd_sc_hd__dfxtp_1 _1883_ (.CLK(clknet_leaf_7_clk),
    .D(_0199_),
    .Q(net51));
 sky130_fd_sc_hd__dfxtp_1 _1884_ (.CLK(clknet_leaf_7_clk),
    .D(_0200_),
    .Q(net52));
 sky130_fd_sc_hd__dfxtp_1 _1885_ (.CLK(clknet_leaf_8_clk),
    .D(net358),
    .Q(net53));
 sky130_fd_sc_hd__dfxtp_1 _1886_ (.CLK(clknet_leaf_8_clk),
    .D(net344),
    .Q(net54));
 sky130_fd_sc_hd__dfxtp_1 _1887_ (.CLK(clknet_leaf_8_clk),
    .D(net373),
    .Q(net56));
 sky130_fd_sc_hd__dfxtp_1 _1888_ (.CLK(clknet_leaf_8_clk),
    .D(net379),
    .Q(net57));
 sky130_fd_sc_hd__dfxtp_1 _1889_ (.CLK(clknet_leaf_21_clk),
    .D(_0205_),
    .Q(net1));
 sky130_fd_sc_hd__dfxtp_1 _1890_ (.CLK(clknet_leaf_21_clk),
    .D(_0206_),
    .Q(net12));
 sky130_fd_sc_hd__dfxtp_1 _1891_ (.CLK(clknet_leaf_21_clk),
    .D(_0207_),
    .Q(net23));
 sky130_fd_sc_hd__dfxtp_1 _1892_ (.CLK(clknet_leaf_21_clk),
    .D(_0208_),
    .Q(net26));
 sky130_fd_sc_hd__dfxtp_1 _1893_ (.CLK(clknet_leaf_21_clk),
    .D(_0209_),
    .Q(net27));
 sky130_fd_sc_hd__dfxtp_1 _1894_ (.CLK(clknet_leaf_21_clk),
    .D(_0210_),
    .Q(net28));
 sky130_fd_sc_hd__dfxtp_1 _1895_ (.CLK(clknet_leaf_21_clk),
    .D(_0211_),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_1 _1896_ (.CLK(clknet_leaf_21_clk),
    .D(_0212_),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_1 _1897_ (.CLK(clknet_leaf_21_clk),
    .D(_0213_),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_1 _1898_ (.CLK(clknet_leaf_21_clk),
    .D(_0214_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_2 _1899_ (.CLK(clknet_leaf_0_clk),
    .D(net211),
    .Q(net2));
 sky130_fd_sc_hd__dfxtp_2 _1900_ (.CLK(clknet_leaf_1_clk),
    .D(net219),
    .Q(net3));
 sky130_fd_sc_hd__dfxtp_2 _1901_ (.CLK(clknet_leaf_1_clk),
    .D(net213),
    .Q(net4));
 sky130_fd_sc_hd__dfxtp_2 _1902_ (.CLK(clknet_leaf_1_clk),
    .D(net221),
    .Q(net5));
 sky130_fd_sc_hd__dfxtp_4 _1903_ (.CLK(clknet_leaf_1_clk),
    .D(net209),
    .Q(net6));
 sky130_fd_sc_hd__dfxtp_4 _1904_ (.CLK(clknet_leaf_1_clk),
    .D(net205),
    .Q(net7));
 sky130_fd_sc_hd__dfxtp_2 _1905_ (.CLK(clknet_leaf_1_clk),
    .D(net207),
    .Q(net8));
 sky130_fd_sc_hd__dfxtp_2 _1906_ (.CLK(clknet_leaf_1_clk),
    .D(net215),
    .Q(net9));
 sky130_fd_sc_hd__dfxtp_4 _1907_ (.CLK(clknet_leaf_1_clk),
    .D(net217),
    .Q(net10));
 sky130_fd_sc_hd__dfxtp_4 _1908_ (.CLK(clknet_leaf_1_clk),
    .D(net203),
    .Q(net11));
 sky130_fd_sc_hd__dfxtp_2 _1909_ (.CLK(clknet_leaf_1_clk),
    .D(net229),
    .Q(net13));
 sky130_fd_sc_hd__dfxtp_2 _1910_ (.CLK(clknet_leaf_1_clk),
    .D(net227),
    .Q(net14));
 sky130_fd_sc_hd__dfxtp_2 _1911_ (.CLK(clknet_leaf_1_clk),
    .D(net225),
    .Q(net15));
 sky130_fd_sc_hd__dfxtp_4 _1912_ (.CLK(clknet_leaf_1_clk),
    .D(net223),
    .Q(net16));
 sky130_fd_sc_hd__dfxtp_2 _1913_ (.CLK(clknet_leaf_6_clk),
    .D(net310),
    .Q(net17));
 sky130_fd_sc_hd__dfxtp_2 _1914_ (.CLK(clknet_leaf_6_clk),
    .D(net312),
    .Q(net18));
 sky130_fd_sc_hd__dfxtp_2 _1915_ (.CLK(clknet_leaf_7_clk),
    .D(_0231_),
    .Q(net19));
 sky130_fd_sc_hd__dfxtp_2 _1916_ (.CLK(clknet_leaf_7_clk),
    .D(_0232_),
    .Q(net20));
 sky130_fd_sc_hd__dfxtp_2 _1917_ (.CLK(clknet_leaf_7_clk),
    .D(_0233_),
    .Q(net21));
 sky130_fd_sc_hd__dfxtp_2 _1918_ (.CLK(clknet_leaf_7_clk),
    .D(_0234_),
    .Q(net22));
 sky130_fd_sc_hd__dfxtp_2 _1919_ (.CLK(clknet_leaf_7_clk),
    .D(_0235_),
    .Q(net24));
 sky130_fd_sc_hd__dfxtp_2 _1920_ (.CLK(clknet_leaf_7_clk),
    .D(_0236_),
    .Q(net25));
 sky130_fd_sc_hd__dfxtp_1 _1921_ (.CLK(clknet_leaf_19_clk),
    .D(_0237_),
    .Q(\forwarding_unit.reg_write_mem ));
 sky130_fd_sc_hd__dfxtp_1 _1922_ (.CLK(clknet_leaf_18_clk),
    .D(_0238_),
    .Q(id_reg_write));
 sky130_fd_sc_hd__dfxtp_1 _1923_ (.CLK(clknet_leaf_19_clk),
    .D(_0239_),
    .Q(\id_alu_src[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1924_ (.CLK(clknet_leaf_20_clk),
    .D(_0240_),
    .Q(\id_ex_rs1_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1925_ (.CLK(clknet_leaf_21_clk),
    .D(_0241_),
    .Q(\id_ex_rs1_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1926_ (.CLK(clknet_leaf_20_clk),
    .D(_0242_),
    .Q(\id_ex_rs1_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1927_ (.CLK(clknet_leaf_21_clk),
    .D(_0243_),
    .Q(\id_ex_rs1_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1928_ (.CLK(clknet_leaf_21_clk),
    .D(_0244_),
    .Q(\id_ex_rs1_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1929_ (.CLK(clknet_leaf_0_clk),
    .D(net265),
    .Q(\id_ex_rs1_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1930_ (.CLK(clknet_leaf_0_clk),
    .D(net261),
    .Q(\id_ex_rs1_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1931_ (.CLK(clknet_leaf_0_clk),
    .D(net259),
    .Q(\id_ex_rs1_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1932_ (.CLK(clknet_leaf_0_clk),
    .D(net285),
    .Q(\id_ex_rs1_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1933_ (.CLK(clknet_leaf_0_clk),
    .D(net299),
    .Q(\id_ex_rs1_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1934_ (.CLK(clknet_leaf_0_clk),
    .D(_0250_),
    .Q(\id_ex_rs1_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1935_ (.CLK(clknet_leaf_0_clk),
    .D(_0251_),
    .Q(\id_ex_rs1_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1936_ (.CLK(clknet_leaf_0_clk),
    .D(_0252_),
    .Q(\id_ex_rs1_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1937_ (.CLK(clknet_leaf_0_clk),
    .D(net360),
    .Q(\id_ex_rs1_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1938_ (.CLK(clknet_leaf_3_clk),
    .D(_0254_),
    .Q(\id_ex_rs1_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1939_ (.CLK(clknet_leaf_3_clk),
    .D(_0255_),
    .Q(\id_ex_rs1_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1940_ (.CLK(clknet_leaf_3_clk),
    .D(_0256_),
    .Q(\id_ex_rs1_data[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1941_ (.CLK(clknet_leaf_0_clk),
    .D(_0257_),
    .Q(\id_ex_rs1_data[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1942_ (.CLK(clknet_leaf_3_clk),
    .D(_0258_),
    .Q(\id_ex_rs1_data[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1943_ (.CLK(clknet_leaf_2_clk),
    .D(_0259_),
    .Q(\id_ex_rs1_data[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1944_ (.CLK(clknet_leaf_0_clk),
    .D(_0260_),
    .Q(\id_ex_rs1_data[20] ));
 sky130_fd_sc_hd__dfxtp_1 _1945_ (.CLK(clknet_leaf_3_clk),
    .D(_0261_),
    .Q(\id_ex_rs1_data[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1946_ (.CLK(clknet_leaf_6_clk),
    .D(_0262_),
    .Q(\id_ex_rs1_data[22] ));
 sky130_fd_sc_hd__dfxtp_1 _1947_ (.CLK(clknet_leaf_5_clk),
    .D(_0263_),
    .Q(\id_ex_rs1_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 _1948_ (.CLK(clknet_leaf_5_clk),
    .D(_0264_),
    .Q(\id_ex_rs1_data[24] ));
 sky130_fd_sc_hd__dfxtp_1 _1949_ (.CLK(clknet_leaf_5_clk),
    .D(_0265_),
    .Q(\id_ex_rs1_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 _1950_ (.CLK(clknet_leaf_5_clk),
    .D(_0266_),
    .Q(\id_ex_rs1_data[26] ));
 sky130_fd_sc_hd__dfxtp_1 _1951_ (.CLK(clknet_leaf_8_clk),
    .D(net340),
    .Q(\id_ex_rs1_data[27] ));
 sky130_fd_sc_hd__dfxtp_1 _1952_ (.CLK(clknet_leaf_8_clk),
    .D(net356),
    .Q(\id_ex_rs1_data[28] ));
 sky130_fd_sc_hd__dfxtp_1 _1953_ (.CLK(clknet_leaf_8_clk),
    .D(net346),
    .Q(\id_ex_rs1_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 _1954_ (.CLK(clknet_leaf_8_clk),
    .D(net354),
    .Q(\id_ex_rs1_data[30] ));
 sky130_fd_sc_hd__dfxtp_1 _1955_ (.CLK(clknet_leaf_8_clk),
    .D(net338),
    .Q(\id_ex_rs1_data[31] ));
 sky130_fd_sc_hd__dfxtp_1 _1956_ (.CLK(clknet_leaf_19_clk),
    .D(_0272_),
    .Q(\id_ex_immediate[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1957_ (.CLK(clknet_leaf_19_clk),
    .D(_0273_),
    .Q(\id_ex_immediate[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1958_ (.CLK(clknet_leaf_19_clk),
    .D(_0274_),
    .Q(\id_ex_immediate[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1959_ (.CLK(clknet_leaf_18_clk),
    .D(_0275_),
    .Q(net103));
 sky130_fd_sc_hd__dfxtp_4 _1960_ (.CLK(clknet_leaf_18_clk),
    .D(_0276_),
    .Q(net97));
 sky130_fd_sc_hd__dfxtp_2 _1961_ (.CLK(clknet_leaf_16_clk),
    .D(_0277_),
    .Q(net100));
 sky130_fd_sc_hd__dfxtp_2 _1962_ (.CLK(clknet_leaf_16_clk),
    .D(_0278_),
    .Q(net99));
 sky130_fd_sc_hd__buf_1 _1989_ (.A(net97),
    .X(net102));
 sky130_fd_sc_hd__buf_1 _1990_ (.A(net99),
    .X(net104));
 sky130_fd_sc_hd__buf_1 _1991_ (.A(net100),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 _1992_ (.A(mem_wb_valid),
    .X(net135));
 sky130_fd_sc_hd__buf_1 _1993_ (.A(ex_mem_valid),
    .X(net136));
 sky130_fd_sc_hd__buf_1 _1994_ (.A(id_ex_valid),
    .X(net137));
 sky130_fd_sc_hd__buf_1 _1995_ (.A(if_id_valid),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(net169),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(net173),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(net174),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(net179),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(net178),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(net183),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(net190),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(net191),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(net193),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(net192),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(net189),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(net187),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(net185),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(net176),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(net179),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(net175),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(net175),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(net180),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(net186),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(net188),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(net182),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(net180),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(net181),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(net177),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(net177),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__inv_8 clkload0 (.A(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload1 (.A(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkinv_4 clkload10 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__inv_8 clkload11 (.A(clknet_leaf_15_clk));
 sky130_fd_sc_hd__inv_8 clkload12 (.A(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkinv_4 clkload13 (.A(clknet_leaf_17_clk));
 sky130_fd_sc_hd__inv_8 clkload14 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkinv_8 clkload2 (.A(clknet_leaf_10_clk));
 sky130_fd_sc_hd__inv_12 clkload3 (.A(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload4 (.A(clknet_leaf_19_clk));
 sky130_fd_sc_hd__inv_6 clkload5 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkinvlp_2 clkload6 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__bufinv_16 clkload7 (.A(clknet_leaf_4_clk));
 sky130_fd_sc_hd__bufinv_16 clkload8 (.A(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkinv_4 clkload9 (.A(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\dmem.address[6] ),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_0220_),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_0174_),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\register_file.write_data[8] ),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_0181_),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(net32),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(_0249_),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\register_file.write_data[0] ),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_0173_),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\register_file.write_data[9] ),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_0182_),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(net47),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\register_file.write_data[16] ),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_0195_),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(net48),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_0196_),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\forwarding_unit.rd_wb[1] ),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_4 hold114 (.A(_0511_),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_0229_),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(net18),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_0230_),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\forwarding_unit.rd_wb[0] ),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_4 hold119 (.A(_0505_),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_0221_),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_0198_),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(net46),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_0194_),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(net49),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_0197_),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(net45),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(_0193_),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\dmem.address[21] ),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(_0022_),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\dmem.address[26] ),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\register_file.write_data[14] ),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(_0027_),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\dmem.address[22] ),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(_0023_),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\dmem.address[23] ),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(_0024_),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(net128),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_0444_),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(_0081_),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\id_ex_rd_addr[0] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(_0076_),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_0219_),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\dmem.address[20] ),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(_0021_),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_4 hold142 (.A(net359),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(_0271_),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(net20),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(_0267_),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\register_file.write_data[29] ),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(_0138_),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(net54),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(_0202_),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\register_file.write_data[10] ),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(net22),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(_0269_),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(net52),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(_0168_),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(net51),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(_0167_),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\register_file.write_data[28] ),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(_0137_),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(net24),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(_0270_),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_0215_),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(net21),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(_0268_),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(net53),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(_0201_),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(net97),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(_0253_),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(net2),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(net3),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(net9),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(net13),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\register_file.write_data[12] ),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(net4),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(net61),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_0147_),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(net62),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(_0148_),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\dmem.address[19] ),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(_0020_),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\register_file.write_data[30] ),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(_0203_),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\dmem.address[17] ),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_0217_),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(_0018_),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\dmem.address[16] ),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(_0017_),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\register_file.write_data[31] ),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(_0204_),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\dmem.address[18] ),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(_0019_),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\dmem.address[14] ),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(net64),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(_0150_),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\register_file.write_data[17] ),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\dmem.address[15] ),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\forwarding_unit.reg_write_wb ),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(net66),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(net67),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(net59),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(_0177_),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(net95),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(net88),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(net89),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(net96),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_0007_),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_0222_),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\id_alu_src[0] ),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(_0597_),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(_0598_),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(_0601_),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(_0626_),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(_0038_),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(net130),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(_0447_),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(_0082_),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(net101),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\register_file.write_data[18] ),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_0502_),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(net56),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(net57),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(net100),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(net19),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\register_file.write_data[26] ),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\ex_mem_alu_result[1] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(ex_mem_valid),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(id_ex_valid),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\dmem.address[11] ),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_0223_),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(net108),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(_0462_),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(_0091_),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\dmem.address[30] ),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(net55),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\dmem.address[10] ),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\dmem.address[25] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\dmem.address[2] ),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\dmem.address[8] ),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\ex_mem_alu_result[0] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\register_file.write_data[11] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\dmem.address[9] ),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(net116),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(_0476_),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(_0099_),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\dmem.address[31] ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\dmem.address[24] ),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(if_id_valid),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\dmem.address[5] ),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\forwarding_unit.reg_write_mem ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(net125),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_0216_),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\dmem.address[28] ),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\dmem.address[3] ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\dmem.address[29] ),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\dmem.address[12] ),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\dmem.address[13] ),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(net93),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\forwarding_unit.rs2_ex[1] ),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(net65),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(net90),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(net76),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\register_file.write_data[13] ),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(net87),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(net94),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(net115),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(_0097_),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(net118),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(_0100_),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(net112),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(_0094_),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(net92),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(net91),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_0218_),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(net121),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(_0103_),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(net107),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(_0461_),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\forwarding_unit.rd_mem[1] ),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(net120),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(_0481_),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(_0102_),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(net114),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(_0471_),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\register_file.write_data[23] ),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(_0096_),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(net111),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(_0466_),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(_0093_),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(net84),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(_0136_),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(net133),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(_0439_),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(_0440_),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(net123),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_0228_),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(_0486_),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(_0105_),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(net27),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(net12),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(net126),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(_0107_),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\register_file.write_data[7] ),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\register_file.write_data[6] ),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(net1),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(net124),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\register_file.write_data[22] ),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(_0106_),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(net26),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(net25),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(net60),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(_0178_),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(net99),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(net132),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(_0451_),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(_0085_),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\register_file.write_data[27] ),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\dmem.address[7] ),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0227_),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\id_ex_rs1_data[26] ),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(_0061_),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(net127),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(net106),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(_0438_),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(net131),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(net23),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(net105),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(_0456_),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(_0087_),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\register_file.write_data[21] ),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(net134),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\id_ex_immediate[0] ),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(_0545_),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(_0547_),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(_0033_),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(id_reg_write),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(net122),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(net119),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(_0101_),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(net110),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0226_),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(_0092_),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(net113),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(_0472_),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(net110),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(net11),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\id_ex_immediate[3] ),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(_0585_),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(_0589_),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(_0036_),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(net15),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\register_file.write_data[20] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(net129),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\id_ex_immediate[1] ),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(_0562_),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(_0563_),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(_0034_),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\id_ex_rs1_data[1] ),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(_0560_),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(_0035_),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(\forwarding_unit.rd_mem[0] ),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(net103),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0225_),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(net17),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\register_file.write_data[29] ),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(net63),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\register_file.write_data[10] ),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(net50),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(net122),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(net119),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\dmem.address[4] ),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_0005_),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net75),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_0128_),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net70),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_0008_),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_0123_),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net72),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_0125_),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net71),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_0124_),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net68),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_0121_),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net73),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_0126_),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net74),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\dmem.address[27] ),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_0127_),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net69),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_0122_),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net79),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_0131_),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net80),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_0132_),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net43),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_0192_),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net40),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0028_),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_0189_),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net39),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_0188_),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net30),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_0247_),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net29),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_0246_),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net38),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_0187_),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net28),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\register_file.write_data[19] ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(_0245_),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net42),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(_0191_),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net41),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_0190_),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net34),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_0183_),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net36),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_0185_),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(net37),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0224_),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_0186_),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(net35),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_0184_),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\register_file.write_data[25] ),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_0134_),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\register_file.write_data[26] ),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_0135_),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\register_file.write_data[24] ),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(_0133_),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(net31),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\register_file.write_data[15] ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_0248_),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(net78),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(_0130_),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(net77),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_0129_),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\register_file.write_data[2] ),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_0175_),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\register_file.write_data[3] ),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_0176_),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\register_file.write_data[1] ),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_1 max_cap1 (.A(_0539_),
    .X(net542));
 sky130_fd_sc_hd__clkbuf_1 max_cap139 (.A(_0623_),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_2 max_cap141 (.A(_0539_),
    .X(net141));
 sky130_fd_sc_hd__buf_1 max_cap142 (.A(net543),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_2 max_length12 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_2 max_length14 (.A(net183),
    .X(net182));
 sky130_fd_sc_hd__buf_1 max_length16 (.A(clknet_1_0__leaf_clk),
    .X(net184));
 sky130_fd_sc_hd__buf_1 max_length18 (.A(net188),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_2 max_length19 (.A(net188),
    .X(net187));
 sky130_fd_sc_hd__buf_1 max_length24 (.A(net193),
    .X(net192));
 sky130_fd_sc_hd__buf_1 max_length26 (.A(net195),
    .X(net194));
 sky130_fd_sc_hd__buf_1 max_length27 (.A(clknet_1_1__leaf_clk),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_2 max_length6 (.A(clknet_0_clk),
    .X(net174));
 sky130_fd_sc_hd__buf_8 output1 (.A(net1),
    .X(debug_reg1[0]));
 sky130_fd_sc_hd__buf_12 output10 (.A(net10),
    .X(debug_reg1[18]));
 sky130_fd_sc_hd__buf_8 output100 (.A(net100),
    .X(instruction_debug[22]));
 sky130_fd_sc_hd__buf_8 output101 (.A(net101),
    .X(instruction_debug[23]));
 sky130_fd_sc_hd__buf_8 output102 (.A(net102),
    .X(instruction_debug[5]));
 sky130_fd_sc_hd__buf_8 output103 (.A(net103),
    .X(instruction_debug[7]));
 sky130_fd_sc_hd__buf_8 output104 (.A(net104),
    .X(instruction_debug[8]));
 sky130_fd_sc_hd__buf_8 output105 (.A(net105),
    .X(pc_current[10]));
 sky130_fd_sc_hd__buf_8 output106 (.A(net106),
    .X(pc_current[11]));
 sky130_fd_sc_hd__buf_8 output107 (.A(net107),
    .X(pc_current[12]));
 sky130_fd_sc_hd__buf_8 output108 (.A(net108),
    .X(pc_current[13]));
 sky130_fd_sc_hd__buf_8 output109 (.A(net109),
    .X(pc_current[14]));
 sky130_fd_sc_hd__buf_12 output11 (.A(net11),
    .X(debug_reg1[19]));
 sky130_fd_sc_hd__buf_8 output110 (.A(net110),
    .X(pc_current[15]));
 sky130_fd_sc_hd__buf_8 output111 (.A(net111),
    .X(pc_current[16]));
 sky130_fd_sc_hd__buf_8 output112 (.A(net112),
    .X(pc_current[17]));
 sky130_fd_sc_hd__buf_8 output113 (.A(net113),
    .X(pc_current[18]));
 sky130_fd_sc_hd__buf_8 output114 (.A(net114),
    .X(pc_current[19]));
 sky130_fd_sc_hd__buf_8 output115 (.A(net115),
    .X(pc_current[20]));
 sky130_fd_sc_hd__buf_8 output116 (.A(net116),
    .X(pc_current[21]));
 sky130_fd_sc_hd__buf_8 output117 (.A(net117),
    .X(pc_current[22]));
 sky130_fd_sc_hd__buf_8 output118 (.A(net118),
    .X(pc_current[23]));
 sky130_fd_sc_hd__buf_8 output119 (.A(net119),
    .X(pc_current[24]));
 sky130_fd_sc_hd__buf_8 output12 (.A(net12),
    .X(debug_reg1[1]));
 sky130_fd_sc_hd__buf_8 output120 (.A(net120),
    .X(pc_current[25]));
 sky130_fd_sc_hd__buf_8 output121 (.A(net121),
    .X(pc_current[26]));
 sky130_fd_sc_hd__buf_8 output122 (.A(net122),
    .X(pc_current[27]));
 sky130_fd_sc_hd__buf_8 output123 (.A(net123),
    .X(pc_current[28]));
 sky130_fd_sc_hd__buf_8 output124 (.A(net124),
    .X(pc_current[29]));
 sky130_fd_sc_hd__buf_8 output125 (.A(net125),
    .X(pc_current[2]));
 sky130_fd_sc_hd__buf_8 output126 (.A(net126),
    .X(pc_current[30]));
 sky130_fd_sc_hd__buf_8 output127 (.A(net127),
    .X(pc_current[31]));
 sky130_fd_sc_hd__buf_8 output128 (.A(net128),
    .X(pc_current[3]));
 sky130_fd_sc_hd__buf_8 output129 (.A(net129),
    .X(pc_current[4]));
 sky130_fd_sc_hd__buf_12 output13 (.A(net13),
    .X(debug_reg1[20]));
 sky130_fd_sc_hd__buf_8 output130 (.A(net130),
    .X(pc_current[5]));
 sky130_fd_sc_hd__buf_8 output131 (.A(net131),
    .X(pc_current[6]));
 sky130_fd_sc_hd__buf_8 output132 (.A(net132),
    .X(pc_current[7]));
 sky130_fd_sc_hd__buf_8 output133 (.A(net133),
    .X(pc_current[8]));
 sky130_fd_sc_hd__buf_8 output134 (.A(net134),
    .X(pc_current[9]));
 sky130_fd_sc_hd__buf_12 output135 (.A(net135),
    .X(pipeline_state[0]));
 sky130_fd_sc_hd__buf_8 output136 (.A(net136),
    .X(pipeline_state[1]));
 sky130_fd_sc_hd__buf_8 output137 (.A(net137),
    .X(pipeline_state[2]));
 sky130_fd_sc_hd__buf_8 output138 (.A(net138),
    .X(pipeline_state[3]));
 sky130_fd_sc_hd__buf_12 output14 (.A(net14),
    .X(debug_reg1[21]));
 sky130_fd_sc_hd__buf_12 output15 (.A(net15),
    .X(debug_reg1[22]));
 sky130_fd_sc_hd__buf_12 output16 (.A(net16),
    .X(debug_reg1[23]));
 sky130_fd_sc_hd__buf_8 output17 (.A(net17),
    .X(debug_reg1[24]));
 sky130_fd_sc_hd__buf_8 output18 (.A(net18),
    .X(debug_reg1[25]));
 sky130_fd_sc_hd__buf_8 output19 (.A(net19),
    .X(debug_reg1[26]));
 sky130_fd_sc_hd__buf_12 output2 (.A(net2),
    .X(debug_reg1[10]));
 sky130_fd_sc_hd__buf_8 output20 (.A(net20),
    .X(debug_reg1[27]));
 sky130_fd_sc_hd__buf_8 output21 (.A(net21),
    .X(debug_reg1[28]));
 sky130_fd_sc_hd__buf_8 output22 (.A(net22),
    .X(debug_reg1[29]));
 sky130_fd_sc_hd__buf_8 output23 (.A(net23),
    .X(debug_reg1[2]));
 sky130_fd_sc_hd__buf_8 output24 (.A(net24),
    .X(debug_reg1[30]));
 sky130_fd_sc_hd__buf_8 output25 (.A(net25),
    .X(debug_reg1[31]));
 sky130_fd_sc_hd__buf_8 output26 (.A(net26),
    .X(debug_reg1[3]));
 sky130_fd_sc_hd__buf_8 output27 (.A(net27),
    .X(debug_reg1[4]));
 sky130_fd_sc_hd__buf_8 output28 (.A(net28),
    .X(debug_reg1[5]));
 sky130_fd_sc_hd__buf_8 output29 (.A(net29),
    .X(debug_reg1[6]));
 sky130_fd_sc_hd__buf_12 output3 (.A(net3),
    .X(debug_reg1[11]));
 sky130_fd_sc_hd__buf_8 output30 (.A(net30),
    .X(debug_reg1[7]));
 sky130_fd_sc_hd__buf_8 output31 (.A(net31),
    .X(debug_reg1[8]));
 sky130_fd_sc_hd__buf_8 output32 (.A(net32),
    .X(debug_reg1[9]));
 sky130_fd_sc_hd__buf_12 output33 (.A(net33),
    .X(debug_reg2[0]));
 sky130_fd_sc_hd__buf_8 output34 (.A(net34),
    .X(debug_reg2[10]));
 sky130_fd_sc_hd__buf_8 output35 (.A(net35),
    .X(debug_reg2[11]));
 sky130_fd_sc_hd__buf_8 output36 (.A(net36),
    .X(debug_reg2[12]));
 sky130_fd_sc_hd__buf_8 output37 (.A(net37),
    .X(debug_reg2[13]));
 sky130_fd_sc_hd__buf_8 output38 (.A(net38),
    .X(debug_reg2[14]));
 sky130_fd_sc_hd__buf_8 output39 (.A(net39),
    .X(debug_reg2[15]));
 sky130_fd_sc_hd__buf_12 output4 (.A(net4),
    .X(debug_reg1[12]));
 sky130_fd_sc_hd__buf_8 output40 (.A(net40),
    .X(debug_reg2[16]));
 sky130_fd_sc_hd__buf_8 output41 (.A(net41),
    .X(debug_reg2[17]));
 sky130_fd_sc_hd__buf_8 output42 (.A(net42),
    .X(debug_reg2[18]));
 sky130_fd_sc_hd__buf_8 output43 (.A(net43),
    .X(debug_reg2[19]));
 sky130_fd_sc_hd__buf_12 output44 (.A(net44),
    .X(debug_reg2[1]));
 sky130_fd_sc_hd__buf_8 output45 (.A(net45),
    .X(debug_reg2[20]));
 sky130_fd_sc_hd__buf_8 output46 (.A(net46),
    .X(debug_reg2[21]));
 sky130_fd_sc_hd__buf_8 output47 (.A(net47),
    .X(debug_reg2[22]));
 sky130_fd_sc_hd__buf_8 output48 (.A(net48),
    .X(debug_reg2[23]));
 sky130_fd_sc_hd__buf_8 output49 (.A(net49),
    .X(debug_reg2[24]));
 sky130_fd_sc_hd__buf_12 output5 (.A(net5),
    .X(debug_reg1[13]));
 sky130_fd_sc_hd__buf_8 output50 (.A(net50),
    .X(debug_reg2[25]));
 sky130_fd_sc_hd__buf_8 output51 (.A(net51),
    .X(debug_reg2[26]));
 sky130_fd_sc_hd__buf_8 output52 (.A(net52),
    .X(debug_reg2[27]));
 sky130_fd_sc_hd__buf_8 output53 (.A(net53),
    .X(debug_reg2[28]));
 sky130_fd_sc_hd__buf_8 output54 (.A(net54),
    .X(debug_reg2[29]));
 sky130_fd_sc_hd__buf_12 output55 (.A(net55),
    .X(debug_reg2[2]));
 sky130_fd_sc_hd__buf_8 output56 (.A(net56),
    .X(debug_reg2[30]));
 sky130_fd_sc_hd__buf_8 output57 (.A(net57),
    .X(debug_reg2[31]));
 sky130_fd_sc_hd__buf_12 output58 (.A(net58),
    .X(debug_reg2[3]));
 sky130_fd_sc_hd__buf_12 output59 (.A(net59),
    .X(debug_reg2[4]));
 sky130_fd_sc_hd__buf_12 output6 (.A(net6),
    .X(debug_reg1[14]));
 sky130_fd_sc_hd__buf_8 output60 (.A(net60),
    .X(debug_reg2[5]));
 sky130_fd_sc_hd__buf_8 output61 (.A(net61),
    .X(debug_reg2[6]));
 sky130_fd_sc_hd__buf_8 output62 (.A(net62),
    .X(debug_reg2[7]));
 sky130_fd_sc_hd__buf_8 output63 (.A(net63),
    .X(debug_reg2[8]));
 sky130_fd_sc_hd__buf_8 output64 (.A(net64),
    .X(debug_reg2[9]));
 sky130_fd_sc_hd__buf_8 output65 (.A(net65),
    .X(debug_reg3[0]));
 sky130_fd_sc_hd__buf_8 output66 (.A(net66),
    .X(debug_reg3[10]));
 sky130_fd_sc_hd__buf_8 output67 (.A(net67),
    .X(debug_reg3[11]));
 sky130_fd_sc_hd__buf_8 output68 (.A(net68),
    .X(debug_reg3[12]));
 sky130_fd_sc_hd__buf_8 output69 (.A(net69),
    .X(debug_reg3[13]));
 sky130_fd_sc_hd__buf_12 output7 (.A(net7),
    .X(debug_reg1[15]));
 sky130_fd_sc_hd__buf_8 output70 (.A(net70),
    .X(debug_reg3[14]));
 sky130_fd_sc_hd__buf_8 output71 (.A(net71),
    .X(debug_reg3[15]));
 sky130_fd_sc_hd__buf_8 output72 (.A(net72),
    .X(debug_reg3[16]));
 sky130_fd_sc_hd__buf_8 output73 (.A(net73),
    .X(debug_reg3[17]));
 sky130_fd_sc_hd__buf_8 output74 (.A(net74),
    .X(debug_reg3[18]));
 sky130_fd_sc_hd__buf_8 output75 (.A(net75),
    .X(debug_reg3[19]));
 sky130_fd_sc_hd__buf_8 output76 (.A(net76),
    .X(debug_reg3[1]));
 sky130_fd_sc_hd__buf_8 output77 (.A(net77),
    .X(debug_reg3[20]));
 sky130_fd_sc_hd__buf_8 output78 (.A(net78),
    .X(debug_reg3[21]));
 sky130_fd_sc_hd__buf_8 output79 (.A(net79),
    .X(debug_reg3[22]));
 sky130_fd_sc_hd__buf_12 output8 (.A(net8),
    .X(debug_reg1[16]));
 sky130_fd_sc_hd__buf_8 output80 (.A(net80),
    .X(debug_reg3[23]));
 sky130_fd_sc_hd__buf_8 output81 (.A(net81),
    .X(debug_reg3[24]));
 sky130_fd_sc_hd__buf_8 output82 (.A(net82),
    .X(debug_reg3[25]));
 sky130_fd_sc_hd__buf_8 output83 (.A(net83),
    .X(debug_reg3[26]));
 sky130_fd_sc_hd__buf_8 output84 (.A(net84),
    .X(debug_reg3[27]));
 sky130_fd_sc_hd__buf_8 output85 (.A(net85),
    .X(debug_reg3[28]));
 sky130_fd_sc_hd__buf_8 output86 (.A(net86),
    .X(debug_reg3[29]));
 sky130_fd_sc_hd__buf_8 output87 (.A(net87),
    .X(debug_reg3[2]));
 sky130_fd_sc_hd__buf_8 output88 (.A(net88),
    .X(debug_reg3[30]));
 sky130_fd_sc_hd__buf_8 output89 (.A(net89),
    .X(debug_reg3[31]));
 sky130_fd_sc_hd__buf_12 output9 (.A(net9),
    .X(debug_reg1[17]));
 sky130_fd_sc_hd__buf_8 output90 (.A(net90),
    .X(debug_reg3[3]));
 sky130_fd_sc_hd__buf_8 output91 (.A(net91),
    .X(debug_reg3[4]));
 sky130_fd_sc_hd__buf_8 output92 (.A(net92),
    .X(debug_reg3[5]));
 sky130_fd_sc_hd__buf_8 output93 (.A(net93),
    .X(debug_reg3[6]));
 sky130_fd_sc_hd__buf_8 output94 (.A(net94),
    .X(debug_reg3[7]));
 sky130_fd_sc_hd__buf_8 output95 (.A(net95),
    .X(debug_reg3[8]));
 sky130_fd_sc_hd__buf_8 output96 (.A(net96),
    .X(debug_reg3[9]));
 sky130_fd_sc_hd__buf_8 output97 (.A(net97),
    .X(instruction_debug[15]));
 sky130_fd_sc_hd__buf_8 output98 (.A(net98),
    .X(instruction_debug[20]));
 sky130_fd_sc_hd__buf_8 output99 (.A(net99),
    .X(instruction_debug[21]));
 sky130_fd_sc_hd__clkbuf_2 wire1 (.A(net170),
    .X(net169));
 sky130_fd_sc_hd__buf_1 wire10 (.A(net182),
    .X(net178));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire11 (.A(net180),
    .X(net179));
 sky130_fd_sc_hd__buf_1 wire13 (.A(net182),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_4 wire140 (.A(net405),
    .X(net140));
 sky130_fd_sc_hd__buf_1 wire15 (.A(clknet_1_0__leaf_clk),
    .X(net183));
 sky130_fd_sc_hd__buf_1 wire17 (.A(net187),
    .X(net185));
 sky130_fd_sc_hd__buf_1 wire2 (.A(net171),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_2 wire20 (.A(clknet_1_1__leaf_clk),
    .X(net188));
 sky130_fd_sc_hd__buf_1 wire21 (.A(net195),
    .X(net189));
 sky130_fd_sc_hd__buf_1 wire22 (.A(net191),
    .X(net190));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire23 (.A(net193),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_2 wire25 (.A(net194),
    .X(net193));
 sky130_fd_sc_hd__buf_1 wire3 (.A(net172),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_1 wire4 (.A(clk),
    .X(net172));
 sky130_fd_sc_hd__buf_1 wire5 (.A(clknet_0_clk),
    .X(net173));
 sky130_fd_sc_hd__buf_1 wire6 (.A(_0536_),
    .X(net543));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire7 (.A(net176),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_2 wire8 (.A(net184),
    .X(net176));
 sky130_fd_sc_hd__dlymetal6s2s_1 wire9 (.A(net178),
    .X(net177));
 assign instruction_debug[0] = net166;
 assign instruction_debug[10] = net147;
 assign instruction_debug[11] = net148;
 assign instruction_debug[12] = net149;
 assign instruction_debug[13] = net150;
 assign instruction_debug[14] = net151;
 assign instruction_debug[16] = net152;
 assign instruction_debug[17] = net153;
 assign instruction_debug[18] = net154;
 assign instruction_debug[19] = net155;
 assign instruction_debug[1] = net167;
 assign instruction_debug[24] = net156;
 assign instruction_debug[25] = net157;
 assign instruction_debug[26] = net158;
 assign instruction_debug[27] = net159;
 assign instruction_debug[28] = net160;
 assign instruction_debug[29] = net161;
 assign instruction_debug[2] = net143;
 assign instruction_debug[30] = net162;
 assign instruction_debug[31] = net163;
 assign instruction_debug[3] = net144;
 assign instruction_debug[4] = net168;
 assign instruction_debug[6] = net145;
 assign instruction_debug[9] = net146;
 assign pc_current[0] = net164;
 assign pc_current[1] = net165;
endmodule
