module CPU_core (clk,
    reset,
    debug_reg1,
    debug_reg2,
    debug_reg3,
    instruction_debug,
    pc_current,
    pipeline_state);
 input clk;
 input reset;
 output [31:0] debug_reg1;
 output [31:0] debug_reg2;
 output [31:0] debug_reg3;
 output [31:0] instruction_debug;
 output [31:0] pc_current;
 output [3:0] pipeline_state;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire \dmem.address[10] ;
 wire \dmem.address[11] ;
 wire \dmem.address[12] ;
 wire \dmem.address[13] ;
 wire \dmem.address[14] ;
 wire \dmem.address[15] ;
 wire \dmem.address[16] ;
 wire \dmem.address[17] ;
 wire \dmem.address[18] ;
 wire \dmem.address[19] ;
 wire \dmem.address[20] ;
 wire \dmem.address[21] ;
 wire \dmem.address[22] ;
 wire \dmem.address[23] ;
 wire \dmem.address[24] ;
 wire \dmem.address[25] ;
 wire \dmem.address[26] ;
 wire \dmem.address[27] ;
 wire \dmem.address[28] ;
 wire \dmem.address[29] ;
 wire \dmem.address[2] ;
 wire \dmem.address[30] ;
 wire \dmem.address[31] ;
 wire \dmem.address[3] ;
 wire \dmem.address[4] ;
 wire \dmem.address[5] ;
 wire \dmem.address[6] ;
 wire \dmem.address[7] ;
 wire \dmem.address[8] ;
 wire \dmem.address[9] ;
 wire \ex_mem_alu_result[0] ;
 wire \ex_mem_alu_result[1] ;
 wire ex_mem_valid;
 wire \forwarding_unit.rd_mem[0] ;
 wire \forwarding_unit.rd_mem[1] ;
 wire \forwarding_unit.rd_wb[0] ;
 wire \forwarding_unit.rd_wb[1] ;
 wire \forwarding_unit.reg_write_mem ;
 wire \forwarding_unit.reg_write_wb ;
 wire \forwarding_unit.rs1_ex[0] ;
 wire \forwarding_unit.rs2_ex[0] ;
 wire \forwarding_unit.rs2_ex[1] ;
 wire \forwarding_unit.rs2_ex[3] ;
 wire \id_alu_src[0] ;
 wire \id_ex_immediate[0] ;
 wire \id_ex_immediate[1] ;
 wire \id_ex_immediate[3] ;
 wire \id_ex_rd_addr[0] ;
 wire \id_ex_rs1_data[0] ;
 wire \id_ex_rs1_data[10] ;
 wire \id_ex_rs1_data[11] ;
 wire \id_ex_rs1_data[12] ;
 wire \id_ex_rs1_data[13] ;
 wire \id_ex_rs1_data[14] ;
 wire \id_ex_rs1_data[15] ;
 wire \id_ex_rs1_data[16] ;
 wire \id_ex_rs1_data[17] ;
 wire \id_ex_rs1_data[18] ;
 wire \id_ex_rs1_data[19] ;
 wire \id_ex_rs1_data[1] ;
 wire \id_ex_rs1_data[20] ;
 wire \id_ex_rs1_data[21] ;
 wire \id_ex_rs1_data[22] ;
 wire \id_ex_rs1_data[23] ;
 wire \id_ex_rs1_data[24] ;
 wire \id_ex_rs1_data[25] ;
 wire \id_ex_rs1_data[26] ;
 wire \id_ex_rs1_data[27] ;
 wire \id_ex_rs1_data[28] ;
 wire \id_ex_rs1_data[29] ;
 wire \id_ex_rs1_data[2] ;
 wire \id_ex_rs1_data[30] ;
 wire \id_ex_rs1_data[31] ;
 wire \id_ex_rs1_data[3] ;
 wire \id_ex_rs1_data[4] ;
 wire \id_ex_rs1_data[5] ;
 wire \id_ex_rs1_data[6] ;
 wire \id_ex_rs1_data[7] ;
 wire \id_ex_rs1_data[8] ;
 wire \id_ex_rs1_data[9] ;
 wire \id_ex_rs2_data[0] ;
 wire \id_ex_rs2_data[10] ;
 wire \id_ex_rs2_data[11] ;
 wire \id_ex_rs2_data[12] ;
 wire \id_ex_rs2_data[13] ;
 wire \id_ex_rs2_data[14] ;
 wire \id_ex_rs2_data[15] ;
 wire \id_ex_rs2_data[16] ;
 wire \id_ex_rs2_data[17] ;
 wire \id_ex_rs2_data[18] ;
 wire \id_ex_rs2_data[19] ;
 wire \id_ex_rs2_data[1] ;
 wire \id_ex_rs2_data[20] ;
 wire \id_ex_rs2_data[21] ;
 wire \id_ex_rs2_data[22] ;
 wire \id_ex_rs2_data[23] ;
 wire \id_ex_rs2_data[24] ;
 wire \id_ex_rs2_data[25] ;
 wire \id_ex_rs2_data[26] ;
 wire \id_ex_rs2_data[27] ;
 wire \id_ex_rs2_data[28] ;
 wire \id_ex_rs2_data[29] ;
 wire \id_ex_rs2_data[2] ;
 wire \id_ex_rs2_data[30] ;
 wire \id_ex_rs2_data[31] ;
 wire \id_ex_rs2_data[3] ;
 wire \id_ex_rs2_data[4] ;
 wire \id_ex_rs2_data[5] ;
 wire \id_ex_rs2_data[6] ;
 wire \id_ex_rs2_data[7] ;
 wire \id_ex_rs2_data[8] ;
 wire \id_ex_rs2_data[9] ;
 wire id_ex_valid;
 wire id_reg_write;
 wire if_id_valid;
 wire mem_wb_valid;
 wire \register_file.write_data[0] ;
 wire \register_file.write_data[10] ;
 wire \register_file.write_data[11] ;
 wire \register_file.write_data[12] ;
 wire \register_file.write_data[13] ;
 wire \register_file.write_data[14] ;
 wire \register_file.write_data[15] ;
 wire \register_file.write_data[16] ;
 wire \register_file.write_data[17] ;
 wire \register_file.write_data[18] ;
 wire \register_file.write_data[19] ;
 wire \register_file.write_data[1] ;
 wire \register_file.write_data[20] ;
 wire \register_file.write_data[21] ;
 wire \register_file.write_data[22] ;
 wire \register_file.write_data[23] ;
 wire \register_file.write_data[24] ;
 wire \register_file.write_data[25] ;
 wire \register_file.write_data[26] ;
 wire \register_file.write_data[27] ;
 wire \register_file.write_data[28] ;
 wire \register_file.write_data[29] ;
 wire \register_file.write_data[2] ;
 wire \register_file.write_data[30] ;
 wire \register_file.write_data[31] ;
 wire \register_file.write_data[3] ;
 wire \register_file.write_data[4] ;
 wire \register_file.write_data[5] ;
 wire \register_file.write_data[6] ;
 wire \register_file.write_data[7] ;
 wire \register_file.write_data[8] ;
 wire \register_file.write_data[9] ;

 sky130_fd_sc_hd__inv_2 _0842_ (.A(reset),
    .Y(_0519_));
 sky130_fd_sc_hd__buf_1 _0843_ (.A(_0519_),
    .X(_0000_));
 sky130_fd_sc_hd__buf_1 _0844_ (.A(_0519_),
    .X(_0520_));
 sky130_fd_sc_hd__and2_2 _0845_ (.A(\ex_mem_alu_result[0] ),
    .B(_0520_),
    .X(_0001_));
 sky130_fd_sc_hd__buf_1 _0846_ (.A(reset),
    .X(_0521_));
 sky130_fd_sc_hd__buf_1 _0847_ (.A(_0521_),
    .X(_0522_));
 sky130_fd_sc_hd__inv_2 _0848_ (.A(\ex_mem_alu_result[1] ),
    .Y(_0523_));
 sky130_fd_sc_hd__nor2_2 _0849_ (.A(_0522_),
    .B(_0523_),
    .Y(_0002_));
 sky130_fd_sc_hd__and2_2 _0850_ (.A(_0000_),
    .B(\dmem.address[2] ),
    .X(_0003_));
 sky130_fd_sc_hd__and2_2 _0851_ (.A(_0000_),
    .B(\dmem.address[3] ),
    .X(_0004_));
 sky130_fd_sc_hd__and2_2 _0852_ (.A(_0000_),
    .B(\dmem.address[4] ),
    .X(_0005_));
 sky130_fd_sc_hd__and2_2 _0853_ (.A(_0000_),
    .B(\dmem.address[5] ),
    .X(_0006_));
 sky130_fd_sc_hd__and2_2 _0854_ (.A(_0000_),
    .B(\dmem.address[6] ),
    .X(_0007_));
 sky130_fd_sc_hd__and2_2 _0855_ (.A(_0000_),
    .B(\dmem.address[7] ),
    .X(_0008_));
 sky130_fd_sc_hd__and2_2 _0856_ (.A(_0000_),
    .B(\dmem.address[8] ),
    .X(_0009_));
 sky130_fd_sc_hd__and2_2 _0857_ (.A(_0000_),
    .B(\dmem.address[9] ),
    .X(_0010_));
 sky130_fd_sc_hd__and2_2 _0858_ (.A(_0000_),
    .B(\dmem.address[10] ),
    .X(_0011_));
 sky130_fd_sc_hd__and2_2 _0859_ (.A(_0000_),
    .B(\dmem.address[11] ),
    .X(_0012_));
 sky130_fd_sc_hd__and2_2 _0860_ (.A(_0000_),
    .B(\dmem.address[12] ),
    .X(_0013_));
 sky130_fd_sc_hd__buf_1 _0861_ (.A(_0519_),
    .X(_0524_));
 sky130_fd_sc_hd__and2_2 _0862_ (.A(_0524_),
    .B(\dmem.address[13] ),
    .X(_0014_));
 sky130_fd_sc_hd__and2_2 _0863_ (.A(_0524_),
    .B(\dmem.address[14] ),
    .X(_0015_));
 sky130_fd_sc_hd__and2_2 _0864_ (.A(_0524_),
    .B(\dmem.address[15] ),
    .X(_0016_));
 sky130_fd_sc_hd__and2_2 _0865_ (.A(_0524_),
    .B(\dmem.address[16] ),
    .X(_0017_));
 sky130_fd_sc_hd__and2_2 _0866_ (.A(_0524_),
    .B(\dmem.address[17] ),
    .X(_0018_));
 sky130_fd_sc_hd__and2_2 _0867_ (.A(_0524_),
    .B(\dmem.address[18] ),
    .X(_0019_));
 sky130_fd_sc_hd__and2_2 _0868_ (.A(_0524_),
    .B(\dmem.address[19] ),
    .X(_0020_));
 sky130_fd_sc_hd__and2_2 _0869_ (.A(_0524_),
    .B(\dmem.address[20] ),
    .X(_0021_));
 sky130_fd_sc_hd__and2_2 _0870_ (.A(_0524_),
    .B(\dmem.address[21] ),
    .X(_0022_));
 sky130_fd_sc_hd__and2_2 _0871_ (.A(_0524_),
    .B(\dmem.address[22] ),
    .X(_0023_));
 sky130_fd_sc_hd__and2_2 _0872_ (.A(_0524_),
    .B(\dmem.address[23] ),
    .X(_0024_));
 sky130_fd_sc_hd__and2_2 _0873_ (.A(_0524_),
    .B(\dmem.address[24] ),
    .X(_0025_));
 sky130_fd_sc_hd__buf_1 _0874_ (.A(_0519_),
    .X(_0525_));
 sky130_fd_sc_hd__and2_2 _0875_ (.A(_0525_),
    .B(\dmem.address[25] ),
    .X(_0026_));
 sky130_fd_sc_hd__and2_2 _0876_ (.A(_0525_),
    .B(\dmem.address[26] ),
    .X(_0027_));
 sky130_fd_sc_hd__and2_2 _0877_ (.A(_0525_),
    .B(\dmem.address[27] ),
    .X(_0028_));
 sky130_fd_sc_hd__and2_2 _0878_ (.A(_0525_),
    .B(\dmem.address[28] ),
    .X(_0029_));
 sky130_fd_sc_hd__and2_2 _0879_ (.A(_0525_),
    .B(\dmem.address[29] ),
    .X(_0030_));
 sky130_fd_sc_hd__and2_2 _0880_ (.A(_0525_),
    .B(\dmem.address[30] ),
    .X(_0031_));
 sky130_fd_sc_hd__and2_2 _0881_ (.A(_0525_),
    .B(\dmem.address[31] ),
    .X(_0032_));
 sky130_fd_sc_hd__o21ai_2 _0882_ (.A1(\forwarding_unit.rd_wb[0] ),
    .A2(\forwarding_unit.rd_wb[1] ),
    .B1(\forwarding_unit.reg_write_wb ),
    .Y(_0526_));
 sky130_fd_sc_hd__or3b_2 _0883_ (.A(\forwarding_unit.rd_wb[1] ),
    .B(_0526_),
    .C_N(\forwarding_unit.rs1_ex[0] ),
    .X(_0527_));
 sky130_fd_sc_hd__buf_1 _0884_ (.A(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__mux2_2 _0885_ (.A0(\register_file.write_data[0] ),
    .A1(\id_ex_rs1_data[0] ),
    .S(_0528_),
    .X(_0529_));
 sky130_fd_sc_hd__o21ai_2 _0886_ (.A1(\forwarding_unit.rd_mem[0] ),
    .A2(\forwarding_unit.rd_mem[1] ),
    .B1(\forwarding_unit.reg_write_mem ),
    .Y(_0530_));
 sky130_fd_sc_hd__or3b_2 _0887_ (.A(_0530_),
    .B(\forwarding_unit.rd_mem[1] ),
    .C_N(\forwarding_unit.rs1_ex[0] ),
    .X(_0531_));
 sky130_fd_sc_hd__buf_1 _0888_ (.A(_0531_),
    .X(_0532_));
 sky130_fd_sc_hd__mux2_2 _0889_ (.A0(\ex_mem_alu_result[0] ),
    .A1(_0529_),
    .S(_0532_),
    .X(_0533_));
 sky130_fd_sc_hd__and2_2 _0890_ (.A(\id_ex_immediate[0] ),
    .B(\id_alu_src[0] ),
    .X(_0534_));
 sky130_fd_sc_hd__o21a_2 _0891_ (.A1(\forwarding_unit.rd_mem[0] ),
    .A2(\forwarding_unit.rd_mem[1] ),
    .B1(\forwarding_unit.reg_write_mem ),
    .X(_0535_));
 sky130_fd_sc_hd__nor4b_2 _0892_ (.A(\forwarding_unit.rd_mem[0] ),
    .B(\forwarding_unit.rs2_ex[3] ),
    .C(\forwarding_unit.rs2_ex[0] ),
    .D_N(\forwarding_unit.rs2_ex[1] ),
    .Y(_0536_));
 sky130_fd_sc_hd__nand2_2 _0893_ (.A(_0535_),
    .B(_0536_),
    .Y(_0537_));
 sky130_fd_sc_hd__o21a_2 _0894_ (.A1(\forwarding_unit.rd_wb[0] ),
    .A2(\forwarding_unit.rd_wb[1] ),
    .B1(\forwarding_unit.reg_write_wb ),
    .X(_0538_));
 sky130_fd_sc_hd__nor4b_2 _0895_ (.A(\forwarding_unit.rd_wb[0] ),
    .B(\forwarding_unit.rs2_ex[3] ),
    .C(\forwarding_unit.rs2_ex[0] ),
    .D_N(\forwarding_unit.rs2_ex[1] ),
    .Y(_0539_));
 sky130_fd_sc_hd__a32o_2 _0896_ (.A1(\register_file.write_data[0] ),
    .A2(_0538_),
    .A3(_0539_),
    .B1(_0535_),
    .B2(_0536_),
    .X(_0540_));
 sky130_fd_sc_hd__or4b_2 _0897_ (.A(\forwarding_unit.rd_wb[0] ),
    .B(\forwarding_unit.rs2_ex[3] ),
    .C(\forwarding_unit.rs2_ex[0] ),
    .D_N(\forwarding_unit.rs2_ex[1] ),
    .X(_0541_));
 sky130_fd_sc_hd__o21a_2 _0898_ (.A1(_0526_),
    .A2(_0541_),
    .B1(\id_ex_rs2_data[0] ),
    .X(_0542_));
 sky130_fd_sc_hd__inv_2 _0899_ (.A(\id_alu_src[0] ),
    .Y(_0543_));
 sky130_fd_sc_hd__o221a_2 _0900_ (.A1(\ex_mem_alu_result[0] ),
    .A2(_0537_),
    .B1(_0540_),
    .B2(_0542_),
    .C1(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__or2_2 _0901_ (.A(_0534_),
    .B(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__or2b_2 _0902_ (.A(_0533_),
    .B_N(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__or2b_2 _0903_ (.A(_0545_),
    .B_N(_0533_),
    .X(_0547_));
 sky130_fd_sc_hd__a21oi_2 _0904_ (.A1(_0546_),
    .A2(_0547_),
    .B1(_0522_),
    .Y(_0033_));
 sky130_fd_sc_hd__or2_2 _0905_ (.A(_0543_),
    .B(\id_ex_immediate[1] ),
    .X(_0548_));
 sky130_fd_sc_hd__or3_2 _0906_ (.A(\register_file.write_data[1] ),
    .B(_0526_),
    .C(_0541_),
    .X(_0549_));
 sky130_fd_sc_hd__a21o_2 _0907_ (.A1(_0538_),
    .A2(_0539_),
    .B1(\id_ex_rs2_data[1] ),
    .X(_0550_));
 sky130_fd_sc_hd__a31o_2 _0908_ (.A1(\ex_mem_alu_result[1] ),
    .A2(_0535_),
    .A3(_0536_),
    .B1(\id_alu_src[0] ),
    .X(_0551_));
 sky130_fd_sc_hd__a31o_2 _0909_ (.A1(_0537_),
    .A2(_0549_),
    .A3(_0550_),
    .B1(_0551_),
    .X(_0552_));
 sky130_fd_sc_hd__a211o_2 _0910_ (.A1(_0548_),
    .A2(_0552_),
    .B1(_0534_),
    .C1(_0544_),
    .X(_0553_));
 sky130_fd_sc_hd__o211ai_2 _0911_ (.A1(_0534_),
    .A2(_0544_),
    .B1(_0548_),
    .C1(_0552_),
    .Y(_0554_));
 sky130_fd_sc_hd__and3b_2 _0912_ (.A_N(\forwarding_unit.rd_mem[1] ),
    .B(\forwarding_unit.rs1_ex[0] ),
    .C(_0535_),
    .X(_0555_));
 sky130_fd_sc_hd__buf_1 _0913_ (.A(_0555_),
    .X(_0556_));
 sky130_fd_sc_hd__nand2_2 _0914_ (.A(\id_ex_rs1_data[1] ),
    .B(_0528_),
    .Y(_0557_));
 sky130_fd_sc_hd__and3b_2 _0915_ (.A_N(\forwarding_unit.rd_wb[1] ),
    .B(_0538_),
    .C(\forwarding_unit.rs1_ex[0] ),
    .X(_0558_));
 sky130_fd_sc_hd__a21oi_2 _0916_ (.A1(\register_file.write_data[1] ),
    .A2(_0558_),
    .B1(_0556_),
    .Y(_0559_));
 sky130_fd_sc_hd__a22o_2 _0917_ (.A1(_0523_),
    .A2(_0556_),
    .B1(_0557_),
    .B2(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__a21oi_2 _0918_ (.A1(_0553_),
    .A2(_0554_),
    .B1(_0560_),
    .Y(_0561_));
 sky130_fd_sc_hd__nand3_2 _0919_ (.A(_0553_),
    .B(_0554_),
    .C(_0560_),
    .Y(_0562_));
 sky130_fd_sc_hd__and2b_2 _0920_ (.A_N(_0561_),
    .B(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__buf_1 _0921_ (.A(_0521_),
    .X(_0564_));
 sky130_fd_sc_hd__a21oi_2 _0922_ (.A1(_0546_),
    .A2(_0563_),
    .B1(_0564_),
    .Y(_0565_));
 sky130_fd_sc_hd__o21a_2 _0923_ (.A1(_0546_),
    .A2(_0563_),
    .B1(_0565_),
    .X(_0034_));
 sky130_fd_sc_hd__nand2_2 _0924_ (.A(_0538_),
    .B(_0539_),
    .Y(_0566_));
 sky130_fd_sc_hd__or4b_2 _0925_ (.A(\forwarding_unit.rd_mem[0] ),
    .B(\forwarding_unit.rs2_ex[3] ),
    .C(\forwarding_unit.rs2_ex[0] ),
    .D_N(\forwarding_unit.rs2_ex[1] ),
    .X(_0567_));
 sky130_fd_sc_hd__nor2_2 _0926_ (.A(_0530_),
    .B(_0567_),
    .Y(_0568_));
 sky130_fd_sc_hd__and3_2 _0927_ (.A(\register_file.write_data[2] ),
    .B(_0538_),
    .C(_0539_),
    .X(_0569_));
 sky130_fd_sc_hd__a211o_2 _0928_ (.A1(\id_ex_rs2_data[2] ),
    .A2(_0566_),
    .B1(_0568_),
    .C1(_0569_),
    .X(_0570_));
 sky130_fd_sc_hd__or2_2 _0929_ (.A(\dmem.address[2] ),
    .B(_0537_),
    .X(_0571_));
 sky130_fd_sc_hd__a31o_2 _0930_ (.A1(_0543_),
    .A2(_0570_),
    .A3(_0571_),
    .B1(_0534_),
    .X(_0572_));
 sky130_fd_sc_hd__xor2_2 _0931_ (.A(_0553_),
    .B(_0572_),
    .X(_0573_));
 sky130_fd_sc_hd__mux2_2 _0932_ (.A0(\register_file.write_data[2] ),
    .A1(\id_ex_rs1_data[2] ),
    .S(_0528_),
    .X(_0574_));
 sky130_fd_sc_hd__mux2_2 _0933_ (.A0(\dmem.address[2] ),
    .A1(_0574_),
    .S(_0532_),
    .X(_0575_));
 sky130_fd_sc_hd__xnor2_2 _0934_ (.A(_0573_),
    .B(_0575_),
    .Y(_0576_));
 sky130_fd_sc_hd__a21o_2 _0935_ (.A1(_0546_),
    .A2(_0562_),
    .B1(_0561_),
    .X(_0577_));
 sky130_fd_sc_hd__a21oi_2 _0936_ (.A1(_0576_),
    .A2(_0577_),
    .B1(_0564_),
    .Y(_0578_));
 sky130_fd_sc_hd__o21a_2 _0937_ (.A1(_0576_),
    .A2(_0577_),
    .B1(_0578_),
    .X(_0035_));
 sky130_fd_sc_hd__a21o_2 _0938_ (.A1(_0538_),
    .A2(_0539_),
    .B1(\id_ex_rs2_data[3] ),
    .X(_0579_));
 sky130_fd_sc_hd__o211a_2 _0939_ (.A1(\register_file.write_data[3] ),
    .A2(_0566_),
    .B1(_0537_),
    .C1(_0579_),
    .X(_0580_));
 sky130_fd_sc_hd__a31o_2 _0940_ (.A1(\dmem.address[3] ),
    .A2(_0535_),
    .A3(_0536_),
    .B1(\id_alu_src[0] ),
    .X(_0581_));
 sky130_fd_sc_hd__o22a_2 _0941_ (.A1(_0543_),
    .A2(\id_ex_immediate[3] ),
    .B1(_0580_),
    .B2(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__or3_2 _0942_ (.A(_0553_),
    .B(_0572_),
    .C(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__buf_1 _0943_ (.A(_0583_),
    .X(_0584_));
 sky130_fd_sc_hd__o21ai_2 _0944_ (.A1(_0553_),
    .A2(_0572_),
    .B1(_0582_),
    .Y(_0585_));
 sky130_fd_sc_hd__nand2_2 _0945_ (.A(_0584_),
    .B(_0585_),
    .Y(_0586_));
 sky130_fd_sc_hd__mux2_2 _0946_ (.A0(\register_file.write_data[3] ),
    .A1(\id_ex_rs1_data[3] ),
    .S(_0528_),
    .X(_0587_));
 sky130_fd_sc_hd__mux2_2 _0947_ (.A0(\dmem.address[3] ),
    .A1(_0587_),
    .S(_0532_),
    .X(_0588_));
 sky130_fd_sc_hd__xnor2_2 _0948_ (.A(_0586_),
    .B(_0588_),
    .Y(_0589_));
 sky130_fd_sc_hd__and2b_2 _0949_ (.A_N(_0573_),
    .B(_0575_),
    .X(_0590_));
 sky130_fd_sc_hd__a21oi_2 _0950_ (.A1(_0576_),
    .A2(_0577_),
    .B1(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__buf_1 _0951_ (.A(_0519_),
    .X(_0592_));
 sky130_fd_sc_hd__o21ai_2 _0952_ (.A1(_0589_),
    .A2(_0591_),
    .B1(_0592_),
    .Y(_0593_));
 sky130_fd_sc_hd__a21oi_2 _0953_ (.A1(_0589_),
    .A2(_0591_),
    .B1(_0593_),
    .Y(_0036_));
 sky130_fd_sc_hd__buf_1 _0954_ (.A(_0568_),
    .X(_0594_));
 sky130_fd_sc_hd__mux2_2 _0955_ (.A0(\register_file.write_data[4] ),
    .A1(\id_ex_rs2_data[4] ),
    .S(_0566_),
    .X(_0595_));
 sky130_fd_sc_hd__or2_2 _0956_ (.A(\dmem.address[4] ),
    .B(_0537_),
    .X(_0596_));
 sky130_fd_sc_hd__o211a_2 _0957_ (.A1(_0594_),
    .A2(_0595_),
    .B1(_0596_),
    .C1(_0543_),
    .X(_0597_));
 sky130_fd_sc_hd__xnor2_2 _0958_ (.A(_0584_),
    .B(_0597_),
    .Y(_0598_));
 sky130_fd_sc_hd__mux2_2 _0959_ (.A0(\register_file.write_data[4] ),
    .A1(\id_ex_rs1_data[4] ),
    .S(_0528_),
    .X(_0599_));
 sky130_fd_sc_hd__mux2_2 _0960_ (.A0(\dmem.address[4] ),
    .A1(_0599_),
    .S(_0532_),
    .X(_0600_));
 sky130_fd_sc_hd__nand2_2 _0961_ (.A(_0598_),
    .B(_0600_),
    .Y(_0601_));
 sky130_fd_sc_hd__or2_2 _0962_ (.A(_0598_),
    .B(_0600_),
    .X(_0602_));
 sky130_fd_sc_hd__nand2_2 _0963_ (.A(_0601_),
    .B(_0602_),
    .Y(_0603_));
 sky130_fd_sc_hd__nand2_2 _0964_ (.A(_0586_),
    .B(_0588_),
    .Y(_0604_));
 sky130_fd_sc_hd__o21a_2 _0965_ (.A1(_0589_),
    .A2(_0591_),
    .B1(_0604_),
    .X(_0605_));
 sky130_fd_sc_hd__or2_2 _0966_ (.A(_0603_),
    .B(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__buf_1 _0967_ (.A(_0521_),
    .X(_0607_));
 sky130_fd_sc_hd__a21oi_2 _0968_ (.A1(_0603_),
    .A2(_0605_),
    .B1(_0607_),
    .Y(_0608_));
 sky130_fd_sc_hd__and2_2 _0969_ (.A(_0606_),
    .B(_0608_),
    .X(_0037_));
 sky130_fd_sc_hd__buf_1 _0970_ (.A(_0566_),
    .X(_0609_));
 sky130_fd_sc_hd__mux2_2 _0971_ (.A0(\register_file.write_data[5] ),
    .A1(\id_ex_rs2_data[5] ),
    .S(_0609_),
    .X(_0610_));
 sky130_fd_sc_hd__buf_1 _0972_ (.A(_0537_),
    .X(_0611_));
 sky130_fd_sc_hd__or2_2 _0973_ (.A(\dmem.address[5] ),
    .B(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__buf_1 _0974_ (.A(_0543_),
    .X(_0613_));
 sky130_fd_sc_hd__o211a_2 _0975_ (.A1(_0594_),
    .A2(_0610_),
    .B1(_0612_),
    .C1(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__or2_2 _0976_ (.A(_0597_),
    .B(_0614_),
    .X(_0615_));
 sky130_fd_sc_hd__nor2_2 _0977_ (.A(_0584_),
    .B(_0615_),
    .Y(_0616_));
 sky130_fd_sc_hd__o21a_2 _0978_ (.A1(_0584_),
    .A2(_0597_),
    .B1(_0614_),
    .X(_0617_));
 sky130_fd_sc_hd__buf_1 _0979_ (.A(_0528_),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_2 _0980_ (.A0(\register_file.write_data[5] ),
    .A1(\id_ex_rs1_data[5] ),
    .S(_0618_),
    .X(_0619_));
 sky130_fd_sc_hd__buf_1 _0981_ (.A(_0532_),
    .X(_0620_));
 sky130_fd_sc_hd__mux2_2 _0982_ (.A0(\dmem.address[5] ),
    .A1(_0619_),
    .S(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__o21ai_2 _0983_ (.A1(_0616_),
    .A2(_0617_),
    .B1(_0621_),
    .Y(_0622_));
 sky130_fd_sc_hd__nor3_2 _0984_ (.A(_0616_),
    .B(_0617_),
    .C(_0621_),
    .Y(_0623_));
 sky130_fd_sc_hd__inv_2 _0985_ (.A(_0623_),
    .Y(_0624_));
 sky130_fd_sc_hd__nand2_2 _0986_ (.A(_0622_),
    .B(_0624_),
    .Y(_0625_));
 sky130_fd_sc_hd__a21oi_2 _0987_ (.A1(_0601_),
    .A2(_0606_),
    .B1(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hd__a31o_2 _0988_ (.A1(_0601_),
    .A2(_0606_),
    .A3(_0625_),
    .B1(_0607_),
    .X(_0627_));
 sky130_fd_sc_hd__nor2_2 _0989_ (.A(_0626_),
    .B(_0627_),
    .Y(_0038_));
 sky130_fd_sc_hd__buf_1 _0990_ (.A(_0519_),
    .X(_0628_));
 sky130_fd_sc_hd__mux2_2 _0991_ (.A0(\register_file.write_data[6] ),
    .A1(\id_ex_rs2_data[6] ),
    .S(_0566_),
    .X(_0629_));
 sky130_fd_sc_hd__or2_2 _0992_ (.A(\dmem.address[6] ),
    .B(_0537_),
    .X(_0630_));
 sky130_fd_sc_hd__o211a_2 _0993_ (.A1(_0594_),
    .A2(_0629_),
    .B1(_0630_),
    .C1(_0543_),
    .X(_0631_));
 sky130_fd_sc_hd__xnor2_2 _0994_ (.A(_0616_),
    .B(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hd__mux2_2 _0995_ (.A0(\register_file.write_data[6] ),
    .A1(\id_ex_rs1_data[6] ),
    .S(_0618_),
    .X(_0633_));
 sky130_fd_sc_hd__mux2_2 _0996_ (.A0(\dmem.address[6] ),
    .A1(_0633_),
    .S(_0620_),
    .X(_0634_));
 sky130_fd_sc_hd__or2b_2 _0997_ (.A(_0632_),
    .B_N(_0634_),
    .X(_0635_));
 sky130_fd_sc_hd__or2b_2 _0998_ (.A(_0634_),
    .B_N(_0632_),
    .X(_0636_));
 sky130_fd_sc_hd__nand2_2 _0999_ (.A(_0635_),
    .B(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__o211a_2 _1000_ (.A1(_0603_),
    .A2(_0605_),
    .B1(_0622_),
    .C1(_0601_),
    .X(_0638_));
 sky130_fd_sc_hd__or2_2 _1001_ (.A(_0623_),
    .B(_0638_),
    .X(_0639_));
 sky130_fd_sc_hd__nand2_2 _1002_ (.A(_0637_),
    .B(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__or2_2 _1003_ (.A(_0637_),
    .B(_0639_),
    .X(_0641_));
 sky130_fd_sc_hd__and3_2 _1004_ (.A(_0628_),
    .B(_0640_),
    .C(_0641_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_2 _1005_ (.A0(\register_file.write_data[7] ),
    .A1(\id_ex_rs2_data[7] ),
    .S(_0566_),
    .X(_0642_));
 sky130_fd_sc_hd__or2_2 _1006_ (.A(\dmem.address[7] ),
    .B(_0537_),
    .X(_0643_));
 sky130_fd_sc_hd__o211a_2 _1007_ (.A1(_0594_),
    .A2(_0642_),
    .B1(_0643_),
    .C1(_0543_),
    .X(_0644_));
 sky130_fd_sc_hd__or2_2 _1008_ (.A(_0631_),
    .B(_0644_),
    .X(_0645_));
 sky130_fd_sc_hd__nor3_2 _1009_ (.A(_0584_),
    .B(_0615_),
    .C(_0645_),
    .Y(_0646_));
 sky130_fd_sc_hd__o31a_2 _1010_ (.A1(_0584_),
    .A2(_0615_),
    .A3(_0631_),
    .B1(_0644_),
    .X(_0647_));
 sky130_fd_sc_hd__or2_2 _1011_ (.A(_0646_),
    .B(_0647_),
    .X(_0648_));
 sky130_fd_sc_hd__mux2_2 _1012_ (.A0(\register_file.write_data[7] ),
    .A1(\id_ex_rs1_data[7] ),
    .S(_0528_),
    .X(_0649_));
 sky130_fd_sc_hd__mux2_2 _1013_ (.A0(\dmem.address[7] ),
    .A1(_0649_),
    .S(_0532_),
    .X(_0650_));
 sky130_fd_sc_hd__nand2_2 _1014_ (.A(_0648_),
    .B(_0650_),
    .Y(_0651_));
 sky130_fd_sc_hd__or3_2 _1015_ (.A(_0646_),
    .B(_0647_),
    .C(_0650_),
    .X(_0652_));
 sky130_fd_sc_hd__nand2_2 _1016_ (.A(_0651_),
    .B(_0652_),
    .Y(_0653_));
 sky130_fd_sc_hd__a21oi_2 _1017_ (.A1(_0635_),
    .A2(_0641_),
    .B1(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__a31o_2 _1018_ (.A1(_0635_),
    .A2(_0641_),
    .A3(_0653_),
    .B1(_0607_),
    .X(_0655_));
 sky130_fd_sc_hd__nor2_2 _1019_ (.A(_0654_),
    .B(_0655_),
    .Y(_0040_));
 sky130_fd_sc_hd__and3b_2 _1020_ (.A_N(_0632_),
    .B(_0634_),
    .C(_0652_),
    .X(_0656_));
 sky130_fd_sc_hd__a21oi_2 _1021_ (.A1(_0648_),
    .A2(_0650_),
    .B1(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__o41a_2 _1022_ (.A1(_0623_),
    .A2(_0637_),
    .A3(_0638_),
    .A4(_0653_),
    .B1(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__or3_2 _1023_ (.A(_0584_),
    .B(_0615_),
    .C(_0645_),
    .X(_0659_));
 sky130_fd_sc_hd__buf_1 _1024_ (.A(_0659_),
    .X(_0660_));
 sky130_fd_sc_hd__and3_2 _1025_ (.A(\register_file.write_data[8] ),
    .B(_0538_),
    .C(_0539_),
    .X(_0661_));
 sky130_fd_sc_hd__o21a_2 _1026_ (.A1(_0526_),
    .A2(_0541_),
    .B1(\id_ex_rs2_data[8] ),
    .X(_0662_));
 sky130_fd_sc_hd__or3_2 _1027_ (.A(\dmem.address[8] ),
    .B(_0530_),
    .C(_0567_),
    .X(_0663_));
 sky130_fd_sc_hd__o311a_2 _1028_ (.A1(_0568_),
    .A2(_0661_),
    .A3(_0662_),
    .B1(_0663_),
    .C1(_0543_),
    .X(_0664_));
 sky130_fd_sc_hd__xnor2_2 _1029_ (.A(_0660_),
    .B(_0664_),
    .Y(_0665_));
 sky130_fd_sc_hd__mux2_2 _1030_ (.A0(\register_file.write_data[8] ),
    .A1(\id_ex_rs1_data[8] ),
    .S(_0618_),
    .X(_0666_));
 sky130_fd_sc_hd__mux2_2 _1031_ (.A0(\dmem.address[8] ),
    .A1(_0666_),
    .S(_0620_),
    .X(_0667_));
 sky130_fd_sc_hd__xnor2_2 _1032_ (.A(_0665_),
    .B(_0667_),
    .Y(_0668_));
 sky130_fd_sc_hd__nand2_2 _1033_ (.A(_0658_),
    .B(_0668_),
    .Y(_0669_));
 sky130_fd_sc_hd__or2_2 _1034_ (.A(_0658_),
    .B(_0668_),
    .X(_0670_));
 sky130_fd_sc_hd__and3_2 _1035_ (.A(_0628_),
    .B(_0669_),
    .C(_0670_),
    .X(_0041_));
 sky130_fd_sc_hd__nand2_2 _1036_ (.A(_0665_),
    .B(_0667_),
    .Y(_0671_));
 sky130_fd_sc_hd__or4_2 _1037_ (.A(_0584_),
    .B(_0615_),
    .C(_0645_),
    .D(_0664_),
    .X(_0672_));
 sky130_fd_sc_hd__and3_2 _1038_ (.A(\register_file.write_data[9] ),
    .B(_0538_),
    .C(_0539_),
    .X(_0673_));
 sky130_fd_sc_hd__o21a_2 _1039_ (.A1(_0526_),
    .A2(_0541_),
    .B1(\id_ex_rs2_data[9] ),
    .X(_0674_));
 sky130_fd_sc_hd__or3_2 _1040_ (.A(\dmem.address[9] ),
    .B(_0530_),
    .C(_0567_),
    .X(_0675_));
 sky130_fd_sc_hd__o311a_2 _1041_ (.A1(_0568_),
    .A2(_0673_),
    .A3(_0674_),
    .B1(_0675_),
    .C1(_0543_),
    .X(_0676_));
 sky130_fd_sc_hd__xnor2_2 _1042_ (.A(_0672_),
    .B(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__mux2_2 _1043_ (.A0(\register_file.write_data[9] ),
    .A1(\id_ex_rs1_data[9] ),
    .S(_0618_),
    .X(_0678_));
 sky130_fd_sc_hd__mux2_2 _1044_ (.A0(\dmem.address[9] ),
    .A1(_0678_),
    .S(_0620_),
    .X(_0679_));
 sky130_fd_sc_hd__xnor2_2 _1045_ (.A(_0677_),
    .B(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__a21oi_2 _1046_ (.A1(_0671_),
    .A2(_0670_),
    .B1(_0680_),
    .Y(_0681_));
 sky130_fd_sc_hd__a31o_2 _1047_ (.A1(_0671_),
    .A2(_0670_),
    .A3(_0680_),
    .B1(_0607_),
    .X(_0682_));
 sky130_fd_sc_hd__nor2_2 _1048_ (.A(_0681_),
    .B(_0682_),
    .Y(_0042_));
 sky130_fd_sc_hd__or2_2 _1049_ (.A(_0664_),
    .B(_0676_),
    .X(_0683_));
 sky130_fd_sc_hd__mux2_2 _1050_ (.A0(\register_file.write_data[10] ),
    .A1(\id_ex_rs2_data[10] ),
    .S(_0609_),
    .X(_0684_));
 sky130_fd_sc_hd__or2_2 _1051_ (.A(\dmem.address[10] ),
    .B(_0611_),
    .X(_0685_));
 sky130_fd_sc_hd__o211a_2 _1052_ (.A1(_0594_),
    .A2(_0684_),
    .B1(_0685_),
    .C1(_0613_),
    .X(_0686_));
 sky130_fd_sc_hd__or2_2 _1053_ (.A(_0683_),
    .B(_0686_),
    .X(_0687_));
 sky130_fd_sc_hd__o21ai_2 _1054_ (.A1(_0660_),
    .A2(_0683_),
    .B1(_0686_),
    .Y(_0688_));
 sky130_fd_sc_hd__o21ai_2 _1055_ (.A1(_0660_),
    .A2(_0687_),
    .B1(_0688_),
    .Y(_0689_));
 sky130_fd_sc_hd__buf_1 _1056_ (.A(_0618_),
    .X(_0690_));
 sky130_fd_sc_hd__mux2_2 _1057_ (.A0(\register_file.write_data[10] ),
    .A1(\id_ex_rs1_data[10] ),
    .S(_0690_),
    .X(_0691_));
 sky130_fd_sc_hd__buf_1 _1058_ (.A(_0620_),
    .X(_0692_));
 sky130_fd_sc_hd__mux2_2 _1059_ (.A0(\dmem.address[10] ),
    .A1(_0691_),
    .S(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__xor2_2 _1060_ (.A(_0689_),
    .B(_0693_),
    .X(_0694_));
 sky130_fd_sc_hd__nor2_2 _1061_ (.A(_0677_),
    .B(_0679_),
    .Y(_0695_));
 sky130_fd_sc_hd__nand2_2 _1062_ (.A(_0677_),
    .B(_0679_),
    .Y(_0696_));
 sky130_fd_sc_hd__o21ai_2 _1063_ (.A1(_0671_),
    .A2(_0695_),
    .B1(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__nor2_2 _1064_ (.A(_0668_),
    .B(_0680_),
    .Y(_0698_));
 sky130_fd_sc_hd__and2b_2 _1065_ (.A_N(_0658_),
    .B(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__or2_2 _1066_ (.A(_0697_),
    .B(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__or2_2 _1067_ (.A(_0694_),
    .B(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__nand2_2 _1068_ (.A(_0694_),
    .B(_0700_),
    .Y(_0702_));
 sky130_fd_sc_hd__and3_2 _1069_ (.A(_0628_),
    .B(_0701_),
    .C(_0702_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_2 _1070_ (.A0(\register_file.write_data[11] ),
    .A1(\id_ex_rs2_data[11] ),
    .S(_0609_),
    .X(_0703_));
 sky130_fd_sc_hd__or2_2 _1071_ (.A(\dmem.address[11] ),
    .B(_0611_),
    .X(_0704_));
 sky130_fd_sc_hd__o211a_2 _1072_ (.A1(_0594_),
    .A2(_0703_),
    .B1(_0704_),
    .C1(_0613_),
    .X(_0705_));
 sky130_fd_sc_hd__or2_2 _1073_ (.A(_0687_),
    .B(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__nor2_2 _1074_ (.A(_0660_),
    .B(_0706_),
    .Y(_0707_));
 sky130_fd_sc_hd__o21a_2 _1075_ (.A1(_0660_),
    .A2(_0687_),
    .B1(_0705_),
    .X(_0708_));
 sky130_fd_sc_hd__mux2_2 _1076_ (.A0(\register_file.write_data[11] ),
    .A1(\id_ex_rs1_data[11] ),
    .S(_0528_),
    .X(_0709_));
 sky130_fd_sc_hd__mux2_2 _1077_ (.A0(\dmem.address[11] ),
    .A1(_0709_),
    .S(_0532_),
    .X(_0710_));
 sky130_fd_sc_hd__o21ai_2 _1078_ (.A1(_0707_),
    .A2(_0708_),
    .B1(_0710_),
    .Y(_0711_));
 sky130_fd_sc_hd__or3_2 _1079_ (.A(_0707_),
    .B(_0708_),
    .C(_0710_),
    .X(_0712_));
 sky130_fd_sc_hd__and2_2 _1080_ (.A(_0711_),
    .B(_0712_),
    .X(_0713_));
 sky130_fd_sc_hd__a21bo_2 _1081_ (.A1(_0689_),
    .A2(_0693_),
    .B1_N(_0702_),
    .X(_0714_));
 sky130_fd_sc_hd__a21o_2 _1082_ (.A1(_0713_),
    .A2(_0714_),
    .B1(_0521_),
    .X(_0715_));
 sky130_fd_sc_hd__o21ba_2 _1083_ (.A1(_0713_),
    .A2(_0714_),
    .B1_N(_0715_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_2 _1084_ (.A0(\register_file.write_data[12] ),
    .A1(\id_ex_rs2_data[12] ),
    .S(_0609_),
    .X(_0716_));
 sky130_fd_sc_hd__o21a_2 _1085_ (.A1(\dmem.address[12] ),
    .A2(_0611_),
    .B1(_0613_),
    .X(_0717_));
 sky130_fd_sc_hd__o21ai_2 _1086_ (.A1(_0594_),
    .A2(_0716_),
    .B1(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hd__or3b_2 _1087_ (.A(_0660_),
    .B(_0706_),
    .C_N(_0718_),
    .X(_0719_));
 sky130_fd_sc_hd__nor2_2 _1088_ (.A(_0687_),
    .B(_0705_),
    .Y(_0720_));
 sky130_fd_sc_hd__a21o_2 _1089_ (.A1(_0646_),
    .A2(_0720_),
    .B1(_0718_),
    .X(_0721_));
 sky130_fd_sc_hd__or2_2 _1090_ (.A(\register_file.write_data[12] ),
    .B(_0618_),
    .X(_0722_));
 sky130_fd_sc_hd__o211a_2 _1091_ (.A1(\id_ex_rs1_data[12] ),
    .A2(_0558_),
    .B1(_0722_),
    .C1(_0620_),
    .X(_0723_));
 sky130_fd_sc_hd__a21oi_2 _1092_ (.A1(\dmem.address[12] ),
    .A2(_0556_),
    .B1(_0723_),
    .Y(_0724_));
 sky130_fd_sc_hd__a21o_2 _1093_ (.A1(_0719_),
    .A2(_0721_),
    .B1(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__nand3_2 _1094_ (.A(_0719_),
    .B(_0721_),
    .C(_0724_),
    .Y(_0726_));
 sky130_fd_sc_hd__nand2_2 _1095_ (.A(_0725_),
    .B(_0726_),
    .Y(_0727_));
 sky130_fd_sc_hd__nand4_2 _1096_ (.A(_0694_),
    .B(_0698_),
    .C(_0711_),
    .D(_0712_),
    .Y(_0728_));
 sky130_fd_sc_hd__and3_2 _1097_ (.A(_0689_),
    .B(_0693_),
    .C(_0712_),
    .X(_0729_));
 sky130_fd_sc_hd__inv_2 _1098_ (.A(_0711_),
    .Y(_0730_));
 sky130_fd_sc_hd__a311oi_2 _1099_ (.A1(_0694_),
    .A2(_0697_),
    .A3(_0712_),
    .B1(_0729_),
    .C1(_0730_),
    .Y(_0731_));
 sky130_fd_sc_hd__o21a_2 _1100_ (.A1(_0658_),
    .A2(_0728_),
    .B1(_0731_),
    .X(_0732_));
 sky130_fd_sc_hd__nand2_2 _1101_ (.A(_0727_),
    .B(_0732_),
    .Y(_0733_));
 sky130_fd_sc_hd__or2_2 _1102_ (.A(_0727_),
    .B(_0732_),
    .X(_0734_));
 sky130_fd_sc_hd__and3_2 _1103_ (.A(_0628_),
    .B(_0733_),
    .C(_0734_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_2 _1104_ (.A0(\register_file.write_data[13] ),
    .A1(\id_ex_rs2_data[13] ),
    .S(_0609_),
    .X(_0735_));
 sky130_fd_sc_hd__o21a_2 _1105_ (.A1(\dmem.address[13] ),
    .A2(_0611_),
    .B1(_0613_),
    .X(_0736_));
 sky130_fd_sc_hd__o21ai_2 _1106_ (.A1(_0594_),
    .A2(_0735_),
    .B1(_0736_),
    .Y(_0737_));
 sky130_fd_sc_hd__nand2_2 _1107_ (.A(_0718_),
    .B(_0737_),
    .Y(_0738_));
 sky130_fd_sc_hd__or3_2 _1108_ (.A(_0660_),
    .B(_0706_),
    .C(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__a31o_2 _1109_ (.A1(_0646_),
    .A2(_0720_),
    .A3(_0718_),
    .B1(_0737_),
    .X(_0740_));
 sky130_fd_sc_hd__or2_2 _1110_ (.A(\register_file.write_data[13] ),
    .B(_0528_),
    .X(_0741_));
 sky130_fd_sc_hd__o211a_2 _1111_ (.A1(\id_ex_rs1_data[13] ),
    .A2(_0558_),
    .B1(_0741_),
    .C1(_0532_),
    .X(_0742_));
 sky130_fd_sc_hd__a21oi_2 _1112_ (.A1(\dmem.address[13] ),
    .A2(_0556_),
    .B1(_0742_),
    .Y(_0743_));
 sky130_fd_sc_hd__and3_2 _1113_ (.A(_0739_),
    .B(_0740_),
    .C(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__a21o_2 _1114_ (.A1(_0739_),
    .A2(_0740_),
    .B1(_0743_),
    .X(_0745_));
 sky130_fd_sc_hd__or2b_2 _1115_ (.A(_0744_),
    .B_N(_0745_),
    .X(_0746_));
 sky130_fd_sc_hd__a21oi_2 _1116_ (.A1(_0725_),
    .A2(_0734_),
    .B1(_0746_),
    .Y(_0747_));
 sky130_fd_sc_hd__a31o_2 _1117_ (.A1(_0725_),
    .A2(_0734_),
    .A3(_0746_),
    .B1(_0607_),
    .X(_0748_));
 sky130_fd_sc_hd__nor2_2 _1118_ (.A(_0747_),
    .B(_0748_),
    .Y(_0046_));
 sky130_fd_sc_hd__mux2_2 _1119_ (.A0(\register_file.write_data[14] ),
    .A1(\id_ex_rs2_data[14] ),
    .S(_0609_),
    .X(_0749_));
 sky130_fd_sc_hd__or2_2 _1120_ (.A(\dmem.address[14] ),
    .B(_0611_),
    .X(_0750_));
 sky130_fd_sc_hd__o211a_2 _1121_ (.A1(_0594_),
    .A2(_0749_),
    .B1(_0750_),
    .C1(_0613_),
    .X(_0751_));
 sky130_fd_sc_hd__or2_2 _1122_ (.A(_0738_),
    .B(_0751_),
    .X(_0752_));
 sky130_fd_sc_hd__or3_2 _1123_ (.A(_0660_),
    .B(_0706_),
    .C(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__a21boi_2 _1124_ (.A1(_0739_),
    .A2(_0751_),
    .B1_N(_0753_),
    .Y(_0754_));
 sky130_fd_sc_hd__mux2_2 _1125_ (.A0(\register_file.write_data[14] ),
    .A1(\id_ex_rs1_data[14] ),
    .S(_0618_),
    .X(_0755_));
 sky130_fd_sc_hd__mux2_2 _1126_ (.A0(\dmem.address[14] ),
    .A1(_0755_),
    .S(_0620_),
    .X(_0756_));
 sky130_fd_sc_hd__xor2_2 _1127_ (.A(_0754_),
    .B(_0756_),
    .X(_0757_));
 sky130_fd_sc_hd__o21a_2 _1128_ (.A1(_0725_),
    .A2(_0744_),
    .B1(_0745_),
    .X(_0758_));
 sky130_fd_sc_hd__o21a_2 _1129_ (.A1(_0734_),
    .A2(_0746_),
    .B1(_0758_),
    .X(_0759_));
 sky130_fd_sc_hd__nand2_2 _1130_ (.A(_0757_),
    .B(_0759_),
    .Y(_0760_));
 sky130_fd_sc_hd__or2_2 _1131_ (.A(_0757_),
    .B(_0759_),
    .X(_0761_));
 sky130_fd_sc_hd__and3_2 _1132_ (.A(_0628_),
    .B(_0760_),
    .C(_0761_),
    .X(_0047_));
 sky130_fd_sc_hd__or2b_2 _1133_ (.A(_0754_),
    .B_N(_0756_),
    .X(_0762_));
 sky130_fd_sc_hd__mux2_2 _1134_ (.A0(\register_file.write_data[15] ),
    .A1(\id_ex_rs2_data[15] ),
    .S(_0609_),
    .X(_0763_));
 sky130_fd_sc_hd__or2_2 _1135_ (.A(\dmem.address[15] ),
    .B(_0611_),
    .X(_0764_));
 sky130_fd_sc_hd__o211a_2 _1136_ (.A1(_0594_),
    .A2(_0763_),
    .B1(_0764_),
    .C1(_0613_),
    .X(_0765_));
 sky130_fd_sc_hd__xnor2_2 _1137_ (.A(_0753_),
    .B(_0765_),
    .Y(_0766_));
 sky130_fd_sc_hd__mux2_2 _1138_ (.A0(\register_file.write_data[15] ),
    .A1(\id_ex_rs1_data[15] ),
    .S(_0618_),
    .X(_0767_));
 sky130_fd_sc_hd__mux2_2 _1139_ (.A0(\dmem.address[15] ),
    .A1(_0767_),
    .S(_0620_),
    .X(_0768_));
 sky130_fd_sc_hd__xnor2_2 _1140_ (.A(_0766_),
    .B(_0768_),
    .Y(_0769_));
 sky130_fd_sc_hd__a21oi_2 _1141_ (.A1(_0762_),
    .A2(_0761_),
    .B1(_0769_),
    .Y(_0770_));
 sky130_fd_sc_hd__a31o_2 _1142_ (.A1(_0762_),
    .A2(_0761_),
    .A3(_0769_),
    .B1(_0607_),
    .X(_0771_));
 sky130_fd_sc_hd__nor2_2 _1143_ (.A(_0770_),
    .B(_0771_),
    .Y(_0048_));
 sky130_fd_sc_hd__or4_2 _1144_ (.A(_0660_),
    .B(_0706_),
    .C(_0752_),
    .D(_0765_),
    .X(_0772_));
 sky130_fd_sc_hd__buf_1 _1145_ (.A(_0772_),
    .X(_0773_));
 sky130_fd_sc_hd__mux2_2 _1146_ (.A0(\register_file.write_data[16] ),
    .A1(\id_ex_rs2_data[16] ),
    .S(_0609_),
    .X(_0774_));
 sky130_fd_sc_hd__or2_2 _1147_ (.A(\dmem.address[16] ),
    .B(_0611_),
    .X(_0775_));
 sky130_fd_sc_hd__o211a_2 _1148_ (.A1(_0594_),
    .A2(_0774_),
    .B1(_0775_),
    .C1(_0613_),
    .X(_0776_));
 sky130_fd_sc_hd__xnor2_2 _1149_ (.A(_0773_),
    .B(_0776_),
    .Y(_0777_));
 sky130_fd_sc_hd__mux2_2 _1150_ (.A0(\register_file.write_data[16] ),
    .A1(\id_ex_rs1_data[16] ),
    .S(_0618_),
    .X(_0778_));
 sky130_fd_sc_hd__mux2_2 _1151_ (.A0(\dmem.address[16] ),
    .A1(_0778_),
    .S(_0620_),
    .X(_0779_));
 sky130_fd_sc_hd__nand2_2 _1152_ (.A(_0777_),
    .B(_0779_),
    .Y(_0780_));
 sky130_fd_sc_hd__or2_2 _1153_ (.A(_0777_),
    .B(_0779_),
    .X(_0781_));
 sky130_fd_sc_hd__nand2_2 _1154_ (.A(_0780_),
    .B(_0781_),
    .Y(_0782_));
 sky130_fd_sc_hd__or4_2 _1155_ (.A(_0727_),
    .B(_0746_),
    .C(_0757_),
    .D(_0769_),
    .X(_0783_));
 sky130_fd_sc_hd__or3_2 _1156_ (.A(_0658_),
    .B(_0728_),
    .C(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__nor2_2 _1157_ (.A(_0766_),
    .B(_0768_),
    .Y(_0785_));
 sky130_fd_sc_hd__nand2_2 _1158_ (.A(_0766_),
    .B(_0768_),
    .Y(_0786_));
 sky130_fd_sc_hd__o21a_2 _1159_ (.A1(_0762_),
    .A2(_0785_),
    .B1(_0786_),
    .X(_0787_));
 sky130_fd_sc_hd__or3_2 _1160_ (.A(_0757_),
    .B(_0758_),
    .C(_0769_),
    .X(_0788_));
 sky130_fd_sc_hd__o211a_2 _1161_ (.A1(_0731_),
    .A2(_0783_),
    .B1(_0787_),
    .C1(_0788_),
    .X(_0789_));
 sky130_fd_sc_hd__and2_2 _1162_ (.A(_0784_),
    .B(_0789_),
    .X(_0790_));
 sky130_fd_sc_hd__nand2_2 _1163_ (.A(_0782_),
    .B(_0790_),
    .Y(_0791_));
 sky130_fd_sc_hd__or2_2 _1164_ (.A(_0782_),
    .B(_0790_),
    .X(_0792_));
 sky130_fd_sc_hd__and3_2 _1165_ (.A(_0628_),
    .B(_0791_),
    .C(_0792_),
    .X(_0049_));
 sky130_fd_sc_hd__and4bb_2 _1166_ (.A_N(_0765_),
    .B_N(_0752_),
    .C(_0720_),
    .D(_0646_),
    .X(_0793_));
 sky130_fd_sc_hd__buf_1 _1167_ (.A(_0594_),
    .X(_0794_));
 sky130_fd_sc_hd__mux2_2 _1168_ (.A0(\register_file.write_data[17] ),
    .A1(\id_ex_rs2_data[17] ),
    .S(_0609_),
    .X(_0795_));
 sky130_fd_sc_hd__or2_2 _1169_ (.A(\dmem.address[17] ),
    .B(_0611_),
    .X(_0796_));
 sky130_fd_sc_hd__o211a_2 _1170_ (.A1(_0794_),
    .A2(_0795_),
    .B1(_0796_),
    .C1(_0613_),
    .X(_0797_));
 sky130_fd_sc_hd__nor2_2 _1171_ (.A(_0776_),
    .B(_0797_),
    .Y(_0798_));
 sky130_fd_sc_hd__nand2_2 _1172_ (.A(_0793_),
    .B(_0798_),
    .Y(_0799_));
 sky130_fd_sc_hd__o21ai_2 _1173_ (.A1(_0773_),
    .A2(_0776_),
    .B1(_0797_),
    .Y(_0800_));
 sky130_fd_sc_hd__or2_2 _1174_ (.A(\register_file.write_data[17] ),
    .B(_0618_),
    .X(_0801_));
 sky130_fd_sc_hd__o211a_2 _1175_ (.A1(\id_ex_rs1_data[17] ),
    .A2(_0558_),
    .B1(_0801_),
    .C1(_0620_),
    .X(_0802_));
 sky130_fd_sc_hd__a21oi_2 _1176_ (.A1(\dmem.address[17] ),
    .A2(_0556_),
    .B1(_0802_),
    .Y(_0803_));
 sky130_fd_sc_hd__and3_2 _1177_ (.A(_0799_),
    .B(_0800_),
    .C(_0803_),
    .X(_0804_));
 sky130_fd_sc_hd__a21o_2 _1178_ (.A1(_0799_),
    .A2(_0800_),
    .B1(_0803_),
    .X(_0805_));
 sky130_fd_sc_hd__or2b_2 _1179_ (.A(_0804_),
    .B_N(_0805_),
    .X(_0806_));
 sky130_fd_sc_hd__a21oi_2 _1180_ (.A1(_0780_),
    .A2(_0792_),
    .B1(_0806_),
    .Y(_0807_));
 sky130_fd_sc_hd__a31o_2 _1181_ (.A1(_0780_),
    .A2(_0792_),
    .A3(_0806_),
    .B1(_0607_),
    .X(_0808_));
 sky130_fd_sc_hd__nor2_2 _1182_ (.A(_0807_),
    .B(_0808_),
    .Y(_0050_));
 sky130_fd_sc_hd__mux2_2 _1183_ (.A0(\register_file.write_data[18] ),
    .A1(\id_ex_rs2_data[18] ),
    .S(_0609_),
    .X(_0809_));
 sky130_fd_sc_hd__mux2_2 _1184_ (.A0(\dmem.address[18] ),
    .A1(_0809_),
    .S(_0611_),
    .X(_0810_));
 sky130_fd_sc_hd__nand2_2 _1185_ (.A(_0613_),
    .B(_0810_),
    .Y(_0811_));
 sky130_fd_sc_hd__nand2_2 _1186_ (.A(_0798_),
    .B(_0811_),
    .Y(_0812_));
 sky130_fd_sc_hd__nor2_2 _1187_ (.A(_0773_),
    .B(_0812_),
    .Y(_0813_));
 sky130_fd_sc_hd__a21oi_2 _1188_ (.A1(_0793_),
    .A2(_0798_),
    .B1(_0811_),
    .Y(_0814_));
 sky130_fd_sc_hd__mux2_2 _1189_ (.A0(\register_file.write_data[18] ),
    .A1(\id_ex_rs1_data[18] ),
    .S(_0618_),
    .X(_0815_));
 sky130_fd_sc_hd__mux2_2 _1190_ (.A0(\dmem.address[18] ),
    .A1(_0815_),
    .S(_0620_),
    .X(_0816_));
 sky130_fd_sc_hd__o21a_2 _1191_ (.A1(_0813_),
    .A2(_0814_),
    .B1(_0816_),
    .X(_0817_));
 sky130_fd_sc_hd__nor3_2 _1192_ (.A(_0813_),
    .B(_0814_),
    .C(_0816_),
    .Y(_0818_));
 sky130_fd_sc_hd__or2_2 _1193_ (.A(_0817_),
    .B(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__o21a_2 _1194_ (.A1(_0780_),
    .A2(_0804_),
    .B1(_0805_),
    .X(_0820_));
 sky130_fd_sc_hd__o31a_2 _1195_ (.A1(_0782_),
    .A2(_0790_),
    .A3(_0806_),
    .B1(_0820_),
    .X(_0821_));
 sky130_fd_sc_hd__o21ai_2 _1196_ (.A1(_0819_),
    .A2(_0821_),
    .B1(_0592_),
    .Y(_0822_));
 sky130_fd_sc_hd__a21oi_2 _1197_ (.A1(_0819_),
    .A2(_0821_),
    .B1(_0822_),
    .Y(_0051_));
 sky130_fd_sc_hd__mux2_2 _1198_ (.A0(\register_file.write_data[19] ),
    .A1(\id_ex_rs2_data[19] ),
    .S(_0609_),
    .X(_0823_));
 sky130_fd_sc_hd__or2_2 _1199_ (.A(\dmem.address[19] ),
    .B(_0611_),
    .X(_0824_));
 sky130_fd_sc_hd__o211a_2 _1200_ (.A1(_0794_),
    .A2(_0823_),
    .B1(_0824_),
    .C1(_0613_),
    .X(_0825_));
 sky130_fd_sc_hd__xor2_2 _1201_ (.A(_0813_),
    .B(_0825_),
    .X(_0826_));
 sky130_fd_sc_hd__mux2_2 _1202_ (.A0(\register_file.write_data[19] ),
    .A1(\id_ex_rs1_data[19] ),
    .S(_0690_),
    .X(_0827_));
 sky130_fd_sc_hd__mux2_2 _1203_ (.A0(\dmem.address[19] ),
    .A1(_0827_),
    .S(_0692_),
    .X(_0828_));
 sky130_fd_sc_hd__xnor2_2 _1204_ (.A(_0826_),
    .B(_0828_),
    .Y(_0829_));
 sky130_fd_sc_hd__o21ba_2 _1205_ (.A1(_0819_),
    .A2(_0821_),
    .B1_N(_0817_),
    .X(_0830_));
 sky130_fd_sc_hd__a21oi_2 _1206_ (.A1(_0829_),
    .A2(_0830_),
    .B1(_0564_),
    .Y(_0831_));
 sky130_fd_sc_hd__o21a_2 _1207_ (.A1(_0829_),
    .A2(_0830_),
    .B1(_0831_),
    .X(_0052_));
 sky130_fd_sc_hd__or2_2 _1208_ (.A(_0812_),
    .B(_0825_),
    .X(_0832_));
 sky130_fd_sc_hd__buf_1 _1209_ (.A(_0609_),
    .X(_0833_));
 sky130_fd_sc_hd__mux2_2 _1210_ (.A0(\register_file.write_data[20] ),
    .A1(\id_ex_rs2_data[20] ),
    .S(_0833_),
    .X(_0834_));
 sky130_fd_sc_hd__buf_1 _1211_ (.A(_0611_),
    .X(_0835_));
 sky130_fd_sc_hd__or2_2 _1212_ (.A(\dmem.address[20] ),
    .B(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__buf_1 _1213_ (.A(_0613_),
    .X(_0837_));
 sky130_fd_sc_hd__o211a_2 _1214_ (.A1(_0794_),
    .A2(_0834_),
    .B1(_0836_),
    .C1(_0837_),
    .X(_0838_));
 sky130_fd_sc_hd__or3_2 _1215_ (.A(_0773_),
    .B(_0832_),
    .C(_0838_),
    .X(_0839_));
 sky130_fd_sc_hd__o21ai_2 _1216_ (.A1(_0773_),
    .A2(_0832_),
    .B1(_0838_),
    .Y(_0840_));
 sky130_fd_sc_hd__or2_2 _1217_ (.A(\register_file.write_data[20] ),
    .B(_0528_),
    .X(_0841_));
 sky130_fd_sc_hd__o211a_2 _1218_ (.A1(\id_ex_rs1_data[20] ),
    .A2(_0558_),
    .B1(_0841_),
    .C1(_0532_),
    .X(_0279_));
 sky130_fd_sc_hd__a21oi_2 _1219_ (.A1(\dmem.address[20] ),
    .A2(_0556_),
    .B1(_0279_),
    .Y(_0280_));
 sky130_fd_sc_hd__a21oi_2 _1220_ (.A1(_0839_),
    .A2(_0840_),
    .B1(_0280_),
    .Y(_0281_));
 sky130_fd_sc_hd__and3_2 _1221_ (.A(_0839_),
    .B(_0840_),
    .C(_0280_),
    .X(_0282_));
 sky130_fd_sc_hd__or2_2 _1222_ (.A(_0281_),
    .B(_0282_),
    .X(_0283_));
 sky130_fd_sc_hd__buf_1 _1223_ (.A(_0283_),
    .X(_0284_));
 sky130_fd_sc_hd__or4_2 _1224_ (.A(_0782_),
    .B(_0806_),
    .C(_0819_),
    .D(_0829_),
    .X(_0285_));
 sky130_fd_sc_hd__a21oi_2 _1225_ (.A1(_0826_),
    .A2(_0828_),
    .B1(_0817_),
    .Y(_0286_));
 sky130_fd_sc_hd__nor2_2 _1226_ (.A(_0826_),
    .B(_0828_),
    .Y(_0287_));
 sky130_fd_sc_hd__o32ai_2 _1227_ (.A1(_0819_),
    .A2(_0820_),
    .A3(_0829_),
    .B1(_0286_),
    .B2(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__o21ba_2 _1228_ (.A1(_0790_),
    .A2(_0285_),
    .B1_N(_0288_),
    .X(_0289_));
 sky130_fd_sc_hd__o21ai_2 _1229_ (.A1(_0284_),
    .A2(_0289_),
    .B1(_0519_),
    .Y(_0290_));
 sky130_fd_sc_hd__a21oi_2 _1230_ (.A1(_0284_),
    .A2(_0289_),
    .B1(_0290_),
    .Y(_0053_));
 sky130_fd_sc_hd__mux2_2 _1231_ (.A0(\register_file.write_data[21] ),
    .A1(\id_ex_rs2_data[21] ),
    .S(_0833_),
    .X(_0291_));
 sky130_fd_sc_hd__or2_2 _1232_ (.A(\dmem.address[21] ),
    .B(_0835_),
    .X(_0292_));
 sky130_fd_sc_hd__o211a_2 _1233_ (.A1(_0794_),
    .A2(_0291_),
    .B1(_0292_),
    .C1(_0837_),
    .X(_0293_));
 sky130_fd_sc_hd__nor2_2 _1234_ (.A(_0838_),
    .B(_0293_),
    .Y(_0294_));
 sky130_fd_sc_hd__nor3b_2 _1235_ (.A(_0773_),
    .B(_0832_),
    .C_N(_0294_),
    .Y(_0295_));
 sky130_fd_sc_hd__o31a_2 _1236_ (.A1(_0773_),
    .A2(_0832_),
    .A3(_0838_),
    .B1(_0293_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_2 _1237_ (.A0(\register_file.write_data[21] ),
    .A1(\id_ex_rs1_data[21] ),
    .S(_0618_),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_2 _1238_ (.A0(\dmem.address[21] ),
    .A1(_0297_),
    .S(_0620_),
    .X(_0298_));
 sky130_fd_sc_hd__o21a_2 _1239_ (.A1(_0295_),
    .A2(_0296_),
    .B1(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__or3_2 _1240_ (.A(_0295_),
    .B(_0296_),
    .C(_0298_),
    .X(_0300_));
 sky130_fd_sc_hd__nand2b_2 _1241_ (.A_N(_0299_),
    .B(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__o21ba_2 _1242_ (.A1(_0284_),
    .A2(_0289_),
    .B1_N(_0281_),
    .X(_0302_));
 sky130_fd_sc_hd__xnor2_2 _1243_ (.A(_0301_),
    .B(_0302_),
    .Y(_0303_));
 sky130_fd_sc_hd__nor2_2 _1244_ (.A(_0522_),
    .B(_0303_),
    .Y(_0054_));
 sky130_fd_sc_hd__mux2_2 _1245_ (.A0(\register_file.write_data[22] ),
    .A1(\id_ex_rs2_data[22] ),
    .S(_0833_),
    .X(_0304_));
 sky130_fd_sc_hd__or2_2 _1246_ (.A(\dmem.address[22] ),
    .B(_0835_),
    .X(_0305_));
 sky130_fd_sc_hd__o211a_2 _1247_ (.A1(_0794_),
    .A2(_0304_),
    .B1(_0305_),
    .C1(_0837_),
    .X(_0306_));
 sky130_fd_sc_hd__xor2_2 _1248_ (.A(_0295_),
    .B(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_2 _1249_ (.A0(\register_file.write_data[22] ),
    .A1(\id_ex_rs1_data[22] ),
    .S(_0690_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_2 _1250_ (.A0(\dmem.address[22] ),
    .A1(_0308_),
    .S(_0692_),
    .X(_0309_));
 sky130_fd_sc_hd__nand2_2 _1251_ (.A(_0307_),
    .B(_0309_),
    .Y(_0310_));
 sky130_fd_sc_hd__or2_2 _1252_ (.A(_0307_),
    .B(_0309_),
    .X(_0311_));
 sky130_fd_sc_hd__and2_2 _1253_ (.A(_0310_),
    .B(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__a21o_2 _1254_ (.A1(_0281_),
    .A2(_0300_),
    .B1(_0299_),
    .X(_0313_));
 sky130_fd_sc_hd__nor3_2 _1255_ (.A(_0284_),
    .B(_0289_),
    .C(_0301_),
    .Y(_0314_));
 sky130_fd_sc_hd__or3_2 _1256_ (.A(_0312_),
    .B(_0313_),
    .C(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__o21ai_2 _1257_ (.A1(_0313_),
    .A2(_0314_),
    .B1(_0312_),
    .Y(_0316_));
 sky130_fd_sc_hd__and3_2 _1258_ (.A(_0628_),
    .B(_0315_),
    .C(_0316_),
    .X(_0055_));
 sky130_fd_sc_hd__or4b_2 _1259_ (.A(_0773_),
    .B(_0832_),
    .C(_0306_),
    .D_N(_0294_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_2 _1260_ (.A0(\register_file.write_data[23] ),
    .A1(\id_ex_rs2_data[23] ),
    .S(_0833_),
    .X(_0318_));
 sky130_fd_sc_hd__or2_2 _1261_ (.A(\dmem.address[23] ),
    .B(_0835_),
    .X(_0319_));
 sky130_fd_sc_hd__o211a_2 _1262_ (.A1(_0794_),
    .A2(_0318_),
    .B1(_0319_),
    .C1(_0837_),
    .X(_0320_));
 sky130_fd_sc_hd__xnor2_2 _1263_ (.A(_0317_),
    .B(_0320_),
    .Y(_0321_));
 sky130_fd_sc_hd__mux2_2 _1264_ (.A0(\register_file.write_data[23] ),
    .A1(\id_ex_rs1_data[23] ),
    .S(_0690_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_2 _1265_ (.A0(\dmem.address[23] ),
    .A1(_0322_),
    .S(_0692_),
    .X(_0323_));
 sky130_fd_sc_hd__xnor2_2 _1266_ (.A(_0321_),
    .B(_0323_),
    .Y(_0324_));
 sky130_fd_sc_hd__a21oi_2 _1267_ (.A1(_0310_),
    .A2(_0316_),
    .B1(_0324_),
    .Y(_0325_));
 sky130_fd_sc_hd__a31o_2 _1268_ (.A1(_0310_),
    .A2(_0316_),
    .A3(_0324_),
    .B1(_0607_),
    .X(_0326_));
 sky130_fd_sc_hd__nor2_2 _1269_ (.A(_0325_),
    .B(_0326_),
    .Y(_0056_));
 sky130_fd_sc_hd__xnor2_2 _1270_ (.A(_0307_),
    .B(_0309_),
    .Y(_0327_));
 sky130_fd_sc_hd__or4_2 _1271_ (.A(_0284_),
    .B(_0301_),
    .C(_0327_),
    .D(_0324_),
    .X(_0328_));
 sky130_fd_sc_hd__a211o_2 _1272_ (.A1(_0784_),
    .A2(_0789_),
    .B1(_0285_),
    .C1(_0328_),
    .X(_0329_));
 sky130_fd_sc_hd__nor2_2 _1273_ (.A(_0327_),
    .B(_0324_),
    .Y(_0330_));
 sky130_fd_sc_hd__nor4_2 _1274_ (.A(_0284_),
    .B(_0301_),
    .C(_0327_),
    .D(_0324_),
    .Y(_0331_));
 sky130_fd_sc_hd__a22o_2 _1275_ (.A1(_0307_),
    .A2(_0309_),
    .B1(_0321_),
    .B2(_0323_),
    .X(_0332_));
 sky130_fd_sc_hd__o21a_2 _1276_ (.A1(_0321_),
    .A2(_0323_),
    .B1(_0332_),
    .X(_0333_));
 sky130_fd_sc_hd__a221oi_2 _1277_ (.A1(_0313_),
    .A2(_0330_),
    .B1(_0331_),
    .B2(_0288_),
    .C1(_0333_),
    .Y(_0334_));
 sky130_fd_sc_hd__nor2_2 _1278_ (.A(_0317_),
    .B(_0320_),
    .Y(_0335_));
 sky130_fd_sc_hd__mux2_2 _1279_ (.A0(\register_file.write_data[24] ),
    .A1(\id_ex_rs2_data[24] ),
    .S(_0833_),
    .X(_0336_));
 sky130_fd_sc_hd__or2_2 _1280_ (.A(\dmem.address[24] ),
    .B(_0835_),
    .X(_0337_));
 sky130_fd_sc_hd__o211a_2 _1281_ (.A1(_0794_),
    .A2(_0336_),
    .B1(_0337_),
    .C1(_0837_),
    .X(_0338_));
 sky130_fd_sc_hd__xnor2_2 _1282_ (.A(_0335_),
    .B(_0338_),
    .Y(_0339_));
 sky130_fd_sc_hd__mux2_2 _1283_ (.A0(\register_file.write_data[24] ),
    .A1(\id_ex_rs1_data[24] ),
    .S(_0690_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_2 _1284_ (.A0(\dmem.address[24] ),
    .A1(_0340_),
    .S(_0692_),
    .X(_0341_));
 sky130_fd_sc_hd__xor2_2 _1285_ (.A(_0339_),
    .B(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__a31o_2 _1286_ (.A1(_0329_),
    .A2(_0334_),
    .A3(_0342_),
    .B1(_0521_),
    .X(_0343_));
 sky130_fd_sc_hd__a21o_2 _1287_ (.A1(_0329_),
    .A2(_0334_),
    .B1(_0342_),
    .X(_0344_));
 sky130_fd_sc_hd__nor2b_2 _1288_ (.A(_0343_),
    .B_N(_0344_),
    .Y(_0057_));
 sky130_fd_sc_hd__or2b_2 _1289_ (.A(_0339_),
    .B_N(_0341_),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_2 _1290_ (.A0(\register_file.write_data[25] ),
    .A1(\id_ex_rs2_data[25] ),
    .S(_0833_),
    .X(_0346_));
 sky130_fd_sc_hd__or2_2 _1291_ (.A(\dmem.address[25] ),
    .B(_0835_),
    .X(_0347_));
 sky130_fd_sc_hd__o211a_2 _1292_ (.A1(_0794_),
    .A2(_0346_),
    .B1(_0347_),
    .C1(_0837_),
    .X(_0348_));
 sky130_fd_sc_hd__or4_2 _1293_ (.A(_0317_),
    .B(_0320_),
    .C(_0338_),
    .D(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__buf_1 _1294_ (.A(_0349_),
    .X(_0350_));
 sky130_fd_sc_hd__o31ai_2 _1295_ (.A1(_0317_),
    .A2(_0320_),
    .A3(_0338_),
    .B1(_0348_),
    .Y(_0351_));
 sky130_fd_sc_hd__nand2_2 _1296_ (.A(_0350_),
    .B(_0351_),
    .Y(_0352_));
 sky130_fd_sc_hd__mux2_2 _1297_ (.A0(\register_file.write_data[25] ),
    .A1(\id_ex_rs1_data[25] ),
    .S(_0690_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_2 _1298_ (.A0(\dmem.address[25] ),
    .A1(_0353_),
    .S(_0692_),
    .X(_0354_));
 sky130_fd_sc_hd__and2_2 _1299_ (.A(_0352_),
    .B(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__or2_2 _1300_ (.A(_0352_),
    .B(_0354_),
    .X(_0356_));
 sky130_fd_sc_hd__or2b_2 _1301_ (.A(_0355_),
    .B_N(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__a21oi_2 _1302_ (.A1(_0345_),
    .A2(_0344_),
    .B1(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__a31o_2 _1303_ (.A1(_0345_),
    .A2(_0344_),
    .A3(_0357_),
    .B1(_0607_),
    .X(_0359_));
 sky130_fd_sc_hd__nor2_2 _1304_ (.A(_0358_),
    .B(_0359_),
    .Y(_0058_));
 sky130_fd_sc_hd__a211o_2 _1305_ (.A1(_0329_),
    .A2(_0334_),
    .B1(_0342_),
    .C1(_0357_),
    .X(_0360_));
 sky130_fd_sc_hd__and2b_2 _1306_ (.A_N(_0345_),
    .B(_0356_),
    .X(_0361_));
 sky130_fd_sc_hd__nor2_2 _1307_ (.A(_0355_),
    .B(_0361_),
    .Y(_0362_));
 sky130_fd_sc_hd__mux2_2 _1308_ (.A0(\register_file.write_data[26] ),
    .A1(\id_ex_rs2_data[26] ),
    .S(_0833_),
    .X(_0363_));
 sky130_fd_sc_hd__or2_2 _1309_ (.A(\dmem.address[26] ),
    .B(_0835_),
    .X(_0364_));
 sky130_fd_sc_hd__o211a_2 _1310_ (.A1(_0794_),
    .A2(_0363_),
    .B1(_0364_),
    .C1(_0837_),
    .X(_0365_));
 sky130_fd_sc_hd__xnor2_2 _1311_ (.A(_0350_),
    .B(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__mux2_2 _1312_ (.A0(\register_file.write_data[26] ),
    .A1(\id_ex_rs1_data[26] ),
    .S(_0690_),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_2 _1313_ (.A0(\dmem.address[26] ),
    .A1(_0367_),
    .S(_0692_),
    .X(_0368_));
 sky130_fd_sc_hd__and2_2 _1314_ (.A(_0366_),
    .B(_0368_),
    .X(_0369_));
 sky130_fd_sc_hd__or2_2 _1315_ (.A(_0366_),
    .B(_0368_),
    .X(_0370_));
 sky130_fd_sc_hd__or2b_2 _1316_ (.A(_0369_),
    .B_N(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__a21oi_2 _1317_ (.A1(_0360_),
    .A2(_0362_),
    .B1(_0371_),
    .Y(_0372_));
 sky130_fd_sc_hd__a31o_2 _1318_ (.A1(_0371_),
    .A2(_0360_),
    .A3(_0362_),
    .B1(_0607_),
    .X(_0373_));
 sky130_fd_sc_hd__nor2_2 _1319_ (.A(_0372_),
    .B(_0373_),
    .Y(_0059_));
 sky130_fd_sc_hd__mux2_2 _1320_ (.A0(\register_file.write_data[27] ),
    .A1(\id_ex_rs2_data[27] ),
    .S(_0833_),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_2 _1321_ (.A0(\dmem.address[27] ),
    .A1(_0374_),
    .S(_0835_),
    .X(_0375_));
 sky130_fd_sc_hd__nand2_2 _1322_ (.A(_0837_),
    .B(_0375_),
    .Y(_0376_));
 sky130_fd_sc_hd__inv_2 _1323_ (.A(_0376_),
    .Y(_0377_));
 sky130_fd_sc_hd__or3_2 _1324_ (.A(_0350_),
    .B(_0365_),
    .C(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__o21ai_2 _1325_ (.A1(_0350_),
    .A2(_0365_),
    .B1(_0377_),
    .Y(_0379_));
 sky130_fd_sc_hd__mux2_2 _1326_ (.A0(\register_file.write_data[27] ),
    .A1(\id_ex_rs1_data[27] ),
    .S(_0690_),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_2 _1327_ (.A0(\dmem.address[27] ),
    .A1(_0380_),
    .S(_0692_),
    .X(_0381_));
 sky130_fd_sc_hd__inv_2 _1328_ (.A(_0381_),
    .Y(_0382_));
 sky130_fd_sc_hd__a21oi_2 _1329_ (.A1(_0378_),
    .A2(_0379_),
    .B1(_0382_),
    .Y(_0383_));
 sky130_fd_sc_hd__nand3_2 _1330_ (.A(_0378_),
    .B(_0379_),
    .C(_0382_),
    .Y(_0384_));
 sky130_fd_sc_hd__and2b_2 _1331_ (.A_N(_0383_),
    .B(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__or2_2 _1332_ (.A(_0369_),
    .B(_0372_),
    .X(_0386_));
 sky130_fd_sc_hd__a21oi_2 _1333_ (.A1(_0385_),
    .A2(_0386_),
    .B1(_0564_),
    .Y(_0387_));
 sky130_fd_sc_hd__o21a_2 _1334_ (.A1(_0385_),
    .A2(_0386_),
    .B1(_0387_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_2 _1335_ (.A0(\register_file.write_data[28] ),
    .A1(\id_ex_rs2_data[28] ),
    .S(_0833_),
    .X(_0388_));
 sky130_fd_sc_hd__or2_2 _1336_ (.A(\dmem.address[28] ),
    .B(_0835_),
    .X(_0389_));
 sky130_fd_sc_hd__o211a_2 _1337_ (.A1(_0794_),
    .A2(_0388_),
    .B1(_0389_),
    .C1(_0837_),
    .X(_0390_));
 sky130_fd_sc_hd__xnor2_2 _1338_ (.A(_0378_),
    .B(_0390_),
    .Y(_0391_));
 sky130_fd_sc_hd__mux2_2 _1339_ (.A0(\register_file.write_data[28] ),
    .A1(\id_ex_rs1_data[28] ),
    .S(_0690_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_2 _1340_ (.A0(\dmem.address[28] ),
    .A1(_0392_),
    .S(_0692_),
    .X(_0393_));
 sky130_fd_sc_hd__xnor2_2 _1341_ (.A(_0391_),
    .B(_0393_),
    .Y(_0394_));
 sky130_fd_sc_hd__a21oi_2 _1342_ (.A1(_0369_),
    .A2(_0384_),
    .B1(_0383_),
    .Y(_0395_));
 sky130_fd_sc_hd__a21oi_2 _1343_ (.A1(_0370_),
    .A2(_0384_),
    .B1(_0383_),
    .Y(_0396_));
 sky130_fd_sc_hd__a31o_2 _1344_ (.A1(_0360_),
    .A2(_0362_),
    .A3(_0395_),
    .B1(_0396_),
    .X(_0397_));
 sky130_fd_sc_hd__nor2_2 _1345_ (.A(_0394_),
    .B(_0397_),
    .Y(_0398_));
 sky130_fd_sc_hd__or2_2 _1346_ (.A(_0521_),
    .B(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__a21oi_2 _1347_ (.A1(_0394_),
    .A2(_0397_),
    .B1(_0399_),
    .Y(_0061_));
 sky130_fd_sc_hd__and2_2 _1348_ (.A(_0391_),
    .B(_0393_),
    .X(_0400_));
 sky130_fd_sc_hd__or4_2 _1349_ (.A(_0350_),
    .B(_0365_),
    .C(_0377_),
    .D(_0390_),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_2 _1350_ (.A0(\register_file.write_data[29] ),
    .A1(\id_ex_rs2_data[29] ),
    .S(_0833_),
    .X(_0402_));
 sky130_fd_sc_hd__or2_2 _1351_ (.A(\dmem.address[29] ),
    .B(_0835_),
    .X(_0403_));
 sky130_fd_sc_hd__o211a_2 _1352_ (.A1(_0794_),
    .A2(_0402_),
    .B1(_0403_),
    .C1(_0837_),
    .X(_0404_));
 sky130_fd_sc_hd__xnor2_2 _1353_ (.A(_0401_),
    .B(_0404_),
    .Y(_0405_));
 sky130_fd_sc_hd__mux2_2 _1354_ (.A0(\register_file.write_data[29] ),
    .A1(\id_ex_rs1_data[29] ),
    .S(_0690_),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_2 _1355_ (.A0(\dmem.address[29] ),
    .A1(_0406_),
    .S(_0692_),
    .X(_0407_));
 sky130_fd_sc_hd__xnor2_2 _1356_ (.A(_0405_),
    .B(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__nor3b_2 _1357_ (.A(_0400_),
    .B(_0398_),
    .C_N(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__o21ba_2 _1358_ (.A1(_0400_),
    .A2(_0398_),
    .B1_N(_0408_),
    .X(_0410_));
 sky130_fd_sc_hd__nor3_2 _1359_ (.A(_0522_),
    .B(_0409_),
    .C(_0410_),
    .Y(_0062_));
 sky130_fd_sc_hd__buf_1 _1360_ (.A(_0519_),
    .X(_0411_));
 sky130_fd_sc_hd__nand2_2 _1361_ (.A(_0405_),
    .B(_0407_),
    .Y(_0412_));
 sky130_fd_sc_hd__nor2_2 _1362_ (.A(_0401_),
    .B(_0404_),
    .Y(_0413_));
 sky130_fd_sc_hd__mux2_2 _1363_ (.A0(\register_file.write_data[30] ),
    .A1(\id_ex_rs2_data[30] ),
    .S(_0833_),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_2 _1364_ (.A0(\dmem.address[30] ),
    .A1(_0414_),
    .S(_0835_),
    .X(_0415_));
 sky130_fd_sc_hd__nand2_2 _1365_ (.A(_0837_),
    .B(_0415_),
    .Y(_0416_));
 sky130_fd_sc_hd__xor2_2 _1366_ (.A(_0413_),
    .B(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_2 _1367_ (.A0(\register_file.write_data[30] ),
    .A1(\id_ex_rs1_data[30] ),
    .S(_0690_),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_2 _1368_ (.A0(\dmem.address[30] ),
    .A1(_0418_),
    .S(_0692_),
    .X(_0419_));
 sky130_fd_sc_hd__or2b_2 _1369_ (.A(_0417_),
    .B_N(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__or2b_2 _1370_ (.A(_0419_),
    .B_N(_0417_),
    .X(_0421_));
 sky130_fd_sc_hd__nand2_2 _1371_ (.A(_0420_),
    .B(_0421_),
    .Y(_0422_));
 sky130_fd_sc_hd__or2_2 _1372_ (.A(_0394_),
    .B(_0408_),
    .X(_0423_));
 sky130_fd_sc_hd__a311o_2 _1373_ (.A1(_0360_),
    .A2(_0362_),
    .A3(_0395_),
    .B1(_0396_),
    .C1(_0423_),
    .X(_0424_));
 sky130_fd_sc_hd__o21ai_2 _1374_ (.A1(_0405_),
    .A2(_0407_),
    .B1(_0400_),
    .Y(_0425_));
 sky130_fd_sc_hd__nand4_2 _1375_ (.A(_0412_),
    .B(_0422_),
    .C(_0424_),
    .D(_0425_),
    .Y(_0426_));
 sky130_fd_sc_hd__a31o_2 _1376_ (.A1(_0412_),
    .A2(_0424_),
    .A3(_0425_),
    .B1(_0422_),
    .X(_0427_));
 sky130_fd_sc_hd__and3_2 _1377_ (.A(_0411_),
    .B(_0426_),
    .C(_0427_),
    .X(_0063_));
 sky130_fd_sc_hd__nand2_2 _1378_ (.A(_0413_),
    .B(_0416_),
    .Y(_0428_));
 sky130_fd_sc_hd__mux2_2 _1379_ (.A0(\register_file.write_data[31] ),
    .A1(\id_ex_rs2_data[31] ),
    .S(_0833_),
    .X(_0429_));
 sky130_fd_sc_hd__or2_2 _1380_ (.A(\dmem.address[31] ),
    .B(_0835_),
    .X(_0430_));
 sky130_fd_sc_hd__o211a_2 _1381_ (.A1(_0794_),
    .A2(_0429_),
    .B1(_0430_),
    .C1(_0837_),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_2 _1382_ (.A0(\register_file.write_data[31] ),
    .A1(\id_ex_rs1_data[31] ),
    .S(_0690_),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_2 _1383_ (.A0(\dmem.address[31] ),
    .A1(_0432_),
    .S(_0692_),
    .X(_0433_));
 sky130_fd_sc_hd__xnor2_2 _1384_ (.A(_0431_),
    .B(_0433_),
    .Y(_0434_));
 sky130_fd_sc_hd__xnor2_2 _1385_ (.A(_0428_),
    .B(_0434_),
    .Y(_0435_));
 sky130_fd_sc_hd__a21oi_2 _1386_ (.A1(_0420_),
    .A2(_0427_),
    .B1(_0435_),
    .Y(_0436_));
 sky130_fd_sc_hd__a31o_2 _1387_ (.A1(_0420_),
    .A2(_0427_),
    .A3(_0435_),
    .B1(_0607_),
    .X(_0437_));
 sky130_fd_sc_hd__nor2_2 _1388_ (.A(_0436_),
    .B(_0437_),
    .Y(_0064_));
 sky130_fd_sc_hd__and2_2 _1389_ (.A(_0525_),
    .B(ex_mem_valid),
    .X(_0065_));
 sky130_fd_sc_hd__and2_2 _1390_ (.A(_0525_),
    .B(id_ex_valid),
    .X(_0066_));
 sky130_fd_sc_hd__and2_2 _1391_ (.A(\forwarding_unit.rd_mem[0] ),
    .B(_0628_),
    .X(_0067_));
 sky130_fd_sc_hd__and2_2 _1392_ (.A(\forwarding_unit.rd_mem[1] ),
    .B(_0628_),
    .X(_0068_));
 sky130_fd_sc_hd__or3_2 _1393_ (.A(pc_current[10]),
    .B(pc_current[9]),
    .C(pc_current[11]),
    .X(_0438_));
 sky130_fd_sc_hd__or4_2 _1394_ (.A(pc_current[6]),
    .B(pc_current[5]),
    .C(pc_current[8]),
    .D(pc_current[7]),
    .X(_0439_));
 sky130_fd_sc_hd__or4_2 _1395_ (.A(reset),
    .B(pc_current[4]),
    .C(_0438_),
    .D(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__nor3b_2 _1396_ (.A(_0440_),
    .B(pc_current[3]),
    .C_N(pc_current[2]),
    .Y(_0069_));
 sky130_fd_sc_hd__buf_1 _1397_ (.A(instruction_debug[15]),
    .X(_0441_));
 sky130_fd_sc_hd__and2_2 _1398_ (.A(_0441_),
    .B(_0628_),
    .X(_0070_));
 sky130_fd_sc_hd__and2_2 _1399_ (.A(_0519_),
    .B(instruction_debug[21]),
    .X(_0071_));
 sky130_fd_sc_hd__and2_2 _1400_ (.A(_0525_),
    .B(instruction_debug[22]),
    .X(_0072_));
 sky130_fd_sc_hd__and2_2 _1401_ (.A(_0525_),
    .B(instruction_debug[23]),
    .X(_0073_));
 sky130_fd_sc_hd__and2_2 _1402_ (.A(_0525_),
    .B(instruction_debug[7]),
    .X(_0074_));
 sky130_fd_sc_hd__buf_1 _1403_ (.A(_0519_),
    .X(_0442_));
 sky130_fd_sc_hd__and2_2 _1404_ (.A(_0442_),
    .B(if_id_valid),
    .X(_0075_));
 sky130_fd_sc_hd__and2_2 _1405_ (.A(_0442_),
    .B(\id_ex_rd_addr[0] ),
    .X(_0076_));
 sky130_fd_sc_hd__and2_2 _1406_ (.A(\forwarding_unit.rs2_ex[1] ),
    .B(_0628_),
    .X(_0077_));
 sky130_fd_sc_hd__and2_2 _1407_ (.A(\forwarding_unit.reg_write_mem ),
    .B(_0628_),
    .X(_0078_));
 sky130_fd_sc_hd__nor2_2 _1408_ (.A(_0522_),
    .B(pc_current[2]),
    .Y(_0079_));
 sky130_fd_sc_hd__xnor2_2 _1409_ (.A(pc_current[3]),
    .B(pc_current[2]),
    .Y(_0443_));
 sky130_fd_sc_hd__nor2_2 _1410_ (.A(_0522_),
    .B(_0443_),
    .Y(_0080_));
 sky130_fd_sc_hd__a21oi_2 _1411_ (.A1(pc_current[3]),
    .A2(pc_current[2]),
    .B1(pc_current[4]),
    .Y(_0444_));
 sky130_fd_sc_hd__a31o_2 _1412_ (.A1(pc_current[4]),
    .A2(pc_current[3]),
    .A3(pc_current[2]),
    .B1(_0521_),
    .X(_0445_));
 sky130_fd_sc_hd__nor2_2 _1413_ (.A(_0444_),
    .B(_0445_),
    .Y(_0081_));
 sky130_fd_sc_hd__and4_2 _1414_ (.A(pc_current[4]),
    .B(pc_current[5]),
    .C(pc_current[3]),
    .D(pc_current[2]),
    .X(_0446_));
 sky130_fd_sc_hd__a31o_2 _1415_ (.A1(pc_current[4]),
    .A2(pc_current[3]),
    .A3(pc_current[2]),
    .B1(pc_current[5]),
    .X(_0447_));
 sky130_fd_sc_hd__nand2_2 _1416_ (.A(_0592_),
    .B(_0447_),
    .Y(_0448_));
 sky130_fd_sc_hd__nor2_2 _1417_ (.A(_0446_),
    .B(_0448_),
    .Y(_0082_));
 sky130_fd_sc_hd__a21oi_2 _1418_ (.A1(pc_current[6]),
    .A2(_0446_),
    .B1(_0564_),
    .Y(_0449_));
 sky130_fd_sc_hd__o21a_2 _1419_ (.A1(pc_current[6]),
    .A2(_0446_),
    .B1(_0449_),
    .X(_0083_));
 sky130_fd_sc_hd__a21oi_2 _1420_ (.A1(pc_current[6]),
    .A2(_0446_),
    .B1(pc_current[7]),
    .Y(_0450_));
 sky130_fd_sc_hd__and3_2 _1421_ (.A(pc_current[6]),
    .B(pc_current[7]),
    .C(_0446_),
    .X(_0451_));
 sky130_fd_sc_hd__nor3_2 _1422_ (.A(_0522_),
    .B(_0450_),
    .C(_0451_),
    .Y(_0084_));
 sky130_fd_sc_hd__buf_1 _1423_ (.A(_0521_),
    .X(_0452_));
 sky130_fd_sc_hd__and4_2 _1424_ (.A(pc_current[6]),
    .B(pc_current[8]),
    .C(pc_current[7]),
    .D(_0446_),
    .X(_0453_));
 sky130_fd_sc_hd__nor2_2 _1425_ (.A(_0452_),
    .B(_0453_),
    .Y(_0454_));
 sky130_fd_sc_hd__o21a_2 _1426_ (.A1(pc_current[8]),
    .A2(_0451_),
    .B1(_0454_),
    .X(_0085_));
 sky130_fd_sc_hd__a21oi_2 _1427_ (.A1(pc_current[9]),
    .A2(_0453_),
    .B1(_0564_),
    .Y(_0455_));
 sky130_fd_sc_hd__o21a_2 _1428_ (.A1(pc_current[9]),
    .A2(_0453_),
    .B1(_0455_),
    .X(_0086_));
 sky130_fd_sc_hd__a21oi_2 _1429_ (.A1(pc_current[9]),
    .A2(_0453_),
    .B1(pc_current[10]),
    .Y(_0456_));
 sky130_fd_sc_hd__and3_2 _1430_ (.A(pc_current[10]),
    .B(pc_current[9]),
    .C(_0453_),
    .X(_0457_));
 sky130_fd_sc_hd__nor3_2 _1431_ (.A(_0522_),
    .B(_0456_),
    .C(_0457_),
    .Y(_0087_));
 sky130_fd_sc_hd__and4_2 _1432_ (.A(pc_current[10]),
    .B(pc_current[9]),
    .C(pc_current[11]),
    .D(_0453_),
    .X(_0458_));
 sky130_fd_sc_hd__nor2_2 _1433_ (.A(_0452_),
    .B(_0458_),
    .Y(_0459_));
 sky130_fd_sc_hd__o21a_2 _1434_ (.A1(pc_current[11]),
    .A2(_0457_),
    .B1(_0459_),
    .X(_0088_));
 sky130_fd_sc_hd__a21oi_2 _1435_ (.A1(pc_current[12]),
    .A2(_0458_),
    .B1(_0564_),
    .Y(_0460_));
 sky130_fd_sc_hd__o21a_2 _1436_ (.A1(pc_current[12]),
    .A2(_0458_),
    .B1(_0460_),
    .X(_0089_));
 sky130_fd_sc_hd__a21oi_2 _1437_ (.A1(pc_current[12]),
    .A2(_0458_),
    .B1(pc_current[13]),
    .Y(_0461_));
 sky130_fd_sc_hd__and3_2 _1438_ (.A(pc_current[12]),
    .B(pc_current[13]),
    .C(_0458_),
    .X(_0462_));
 sky130_fd_sc_hd__nor3_2 _1439_ (.A(_0522_),
    .B(_0461_),
    .C(_0462_),
    .Y(_0090_));
 sky130_fd_sc_hd__and2_2 _1440_ (.A(pc_current[14]),
    .B(_0462_),
    .X(_0463_));
 sky130_fd_sc_hd__nor2_2 _1441_ (.A(_0452_),
    .B(_0463_),
    .Y(_0464_));
 sky130_fd_sc_hd__o21a_2 _1442_ (.A1(pc_current[14]),
    .A2(_0462_),
    .B1(_0464_),
    .X(_0091_));
 sky130_fd_sc_hd__a21oi_2 _1443_ (.A1(pc_current[15]),
    .A2(_0463_),
    .B1(_0564_),
    .Y(_0465_));
 sky130_fd_sc_hd__o21a_2 _1444_ (.A1(pc_current[15]),
    .A2(_0463_),
    .B1(_0465_),
    .X(_0092_));
 sky130_fd_sc_hd__a21oi_2 _1445_ (.A1(pc_current[15]),
    .A2(_0463_),
    .B1(pc_current[16]),
    .Y(_0466_));
 sky130_fd_sc_hd__and3_2 _1446_ (.A(pc_current[15]),
    .B(pc_current[16]),
    .C(_0463_),
    .X(_0467_));
 sky130_fd_sc_hd__nor3_2 _1447_ (.A(_0522_),
    .B(_0466_),
    .C(_0467_),
    .Y(_0093_));
 sky130_fd_sc_hd__and2_2 _1448_ (.A(pc_current[17]),
    .B(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__nor2_2 _1449_ (.A(_0452_),
    .B(_0468_),
    .Y(_0469_));
 sky130_fd_sc_hd__o21a_2 _1450_ (.A1(pc_current[17]),
    .A2(_0467_),
    .B1(_0469_),
    .X(_0094_));
 sky130_fd_sc_hd__a21oi_2 _1451_ (.A1(pc_current[18]),
    .A2(_0468_),
    .B1(_0564_),
    .Y(_0470_));
 sky130_fd_sc_hd__o21a_2 _1452_ (.A1(pc_current[18]),
    .A2(_0468_),
    .B1(_0470_),
    .X(_0095_));
 sky130_fd_sc_hd__a21oi_2 _1453_ (.A1(pc_current[18]),
    .A2(_0468_),
    .B1(pc_current[19]),
    .Y(_0471_));
 sky130_fd_sc_hd__and3_2 _1454_ (.A(pc_current[18]),
    .B(pc_current[19]),
    .C(_0468_),
    .X(_0472_));
 sky130_fd_sc_hd__nor3_2 _1455_ (.A(_0522_),
    .B(_0471_),
    .C(_0472_),
    .Y(_0096_));
 sky130_fd_sc_hd__and2_2 _1456_ (.A(pc_current[20]),
    .B(_0472_),
    .X(_0473_));
 sky130_fd_sc_hd__nor2_2 _1457_ (.A(_0452_),
    .B(_0473_),
    .Y(_0474_));
 sky130_fd_sc_hd__o21a_2 _1458_ (.A1(pc_current[20]),
    .A2(_0472_),
    .B1(_0474_),
    .X(_0097_));
 sky130_fd_sc_hd__a21oi_2 _1459_ (.A1(pc_current[21]),
    .A2(_0473_),
    .B1(_0452_),
    .Y(_0475_));
 sky130_fd_sc_hd__o21a_2 _1460_ (.A1(pc_current[21]),
    .A2(_0473_),
    .B1(_0475_),
    .X(_0098_));
 sky130_fd_sc_hd__a21oi_2 _1461_ (.A1(pc_current[21]),
    .A2(_0473_),
    .B1(pc_current[22]),
    .Y(_0476_));
 sky130_fd_sc_hd__and3_2 _1462_ (.A(pc_current[21]),
    .B(pc_current[22]),
    .C(_0473_),
    .X(_0477_));
 sky130_fd_sc_hd__nor3_2 _1463_ (.A(_0564_),
    .B(_0476_),
    .C(_0477_),
    .Y(_0099_));
 sky130_fd_sc_hd__and2_2 _1464_ (.A(pc_current[23]),
    .B(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__nor2_2 _1465_ (.A(_0452_),
    .B(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__o21a_2 _1466_ (.A1(pc_current[23]),
    .A2(_0477_),
    .B1(_0479_),
    .X(_0100_));
 sky130_fd_sc_hd__a21oi_2 _1467_ (.A1(pc_current[24]),
    .A2(_0478_),
    .B1(_0452_),
    .Y(_0480_));
 sky130_fd_sc_hd__o21a_2 _1468_ (.A1(pc_current[24]),
    .A2(_0478_),
    .B1(_0480_),
    .X(_0101_));
 sky130_fd_sc_hd__a21oi_2 _1469_ (.A1(pc_current[24]),
    .A2(_0478_),
    .B1(pc_current[25]),
    .Y(_0481_));
 sky130_fd_sc_hd__and3_2 _1470_ (.A(pc_current[24]),
    .B(pc_current[25]),
    .C(_0478_),
    .X(_0482_));
 sky130_fd_sc_hd__nor3_2 _1471_ (.A(_0564_),
    .B(_0481_),
    .C(_0482_),
    .Y(_0102_));
 sky130_fd_sc_hd__and2_2 _1472_ (.A(pc_current[26]),
    .B(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__nor2_2 _1473_ (.A(_0452_),
    .B(_0483_),
    .Y(_0484_));
 sky130_fd_sc_hd__o21a_2 _1474_ (.A1(pc_current[26]),
    .A2(_0482_),
    .B1(_0484_),
    .X(_0103_));
 sky130_fd_sc_hd__a21oi_2 _1475_ (.A1(pc_current[27]),
    .A2(_0483_),
    .B1(_0452_),
    .Y(_0485_));
 sky130_fd_sc_hd__o21a_2 _1476_ (.A1(pc_current[27]),
    .A2(_0483_),
    .B1(_0485_),
    .X(_0104_));
 sky130_fd_sc_hd__a21oi_2 _1477_ (.A1(pc_current[27]),
    .A2(_0483_),
    .B1(pc_current[28]),
    .Y(_0486_));
 sky130_fd_sc_hd__and3_2 _1478_ (.A(pc_current[27]),
    .B(pc_current[28]),
    .C(_0483_),
    .X(_0487_));
 sky130_fd_sc_hd__nor3_2 _1479_ (.A(_0564_),
    .B(_0486_),
    .C(_0487_),
    .Y(_0105_));
 sky130_fd_sc_hd__and2_2 _1480_ (.A(pc_current[29]),
    .B(_0487_),
    .X(_0488_));
 sky130_fd_sc_hd__nor2_2 _1481_ (.A(_0452_),
    .B(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__o21a_2 _1482_ (.A1(pc_current[29]),
    .A2(_0487_),
    .B1(_0489_),
    .X(_0106_));
 sky130_fd_sc_hd__and3_2 _1483_ (.A(pc_current[29]),
    .B(pc_current[30]),
    .C(_0487_),
    .X(_0490_));
 sky130_fd_sc_hd__nor2_2 _1484_ (.A(_0607_),
    .B(_0490_),
    .Y(_0491_));
 sky130_fd_sc_hd__o21a_2 _1485_ (.A1(pc_current[30]),
    .A2(_0488_),
    .B1(_0491_),
    .X(_0107_));
 sky130_fd_sc_hd__a21oi_2 _1486_ (.A1(pc_current[31]),
    .A2(_0490_),
    .B1(_0452_),
    .Y(_0492_));
 sky130_fd_sc_hd__o21a_2 _1487_ (.A1(pc_current[31]),
    .A2(_0490_),
    .B1(_0492_),
    .X(_0108_));
 sky130_fd_sc_hd__or3b_2 _1488_ (.A(_0526_),
    .B(reset),
    .C_N(mem_wb_valid),
    .X(_0493_));
 sky130_fd_sc_hd__inv_2 _1489_ (.A(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__and3_2 _1490_ (.A(\forwarding_unit.rd_wb[0] ),
    .B(\forwarding_unit.rd_wb[1] ),
    .C(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__buf_1 _1491_ (.A(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__buf_1 _1492_ (.A(_0496_),
    .X(_0497_));
 sky130_fd_sc_hd__nor2_2 _1493_ (.A(_0521_),
    .B(_0496_),
    .Y(_0498_));
 sky130_fd_sc_hd__buf_1 _1494_ (.A(_0498_),
    .X(_0499_));
 sky130_fd_sc_hd__a22o_2 _1495_ (.A1(\register_file.write_data[0] ),
    .A2(_0497_),
    .B1(_0499_),
    .B2(debug_reg3[0]),
    .X(_0109_));
 sky130_fd_sc_hd__a22o_2 _1496_ (.A1(\register_file.write_data[1] ),
    .A2(_0497_),
    .B1(_0499_),
    .B2(debug_reg3[1]),
    .X(_0110_));
 sky130_fd_sc_hd__a22o_2 _1497_ (.A1(\register_file.write_data[2] ),
    .A2(_0497_),
    .B1(_0499_),
    .B2(debug_reg3[2]),
    .X(_0111_));
 sky130_fd_sc_hd__a22o_2 _1498_ (.A1(\register_file.write_data[3] ),
    .A2(_0497_),
    .B1(_0499_),
    .B2(debug_reg3[3]),
    .X(_0112_));
 sky130_fd_sc_hd__a22o_2 _1499_ (.A1(\register_file.write_data[4] ),
    .A2(_0497_),
    .B1(_0499_),
    .B2(debug_reg3[4]),
    .X(_0113_));
 sky130_fd_sc_hd__a22o_2 _1500_ (.A1(\register_file.write_data[5] ),
    .A2(_0497_),
    .B1(_0499_),
    .B2(debug_reg3[5]),
    .X(_0114_));
 sky130_fd_sc_hd__a22o_2 _1501_ (.A1(\register_file.write_data[6] ),
    .A2(_0497_),
    .B1(_0499_),
    .B2(debug_reg3[6]),
    .X(_0115_));
 sky130_fd_sc_hd__a22o_2 _1502_ (.A1(\register_file.write_data[7] ),
    .A2(_0497_),
    .B1(_0499_),
    .B2(debug_reg3[7]),
    .X(_0116_));
 sky130_fd_sc_hd__a22o_2 _1503_ (.A1(\register_file.write_data[8] ),
    .A2(_0497_),
    .B1(_0499_),
    .B2(debug_reg3[8]),
    .X(_0117_));
 sky130_fd_sc_hd__a22o_2 _1504_ (.A1(\register_file.write_data[9] ),
    .A2(_0497_),
    .B1(_0499_),
    .B2(debug_reg3[9]),
    .X(_0118_));
 sky130_fd_sc_hd__a22o_2 _1505_ (.A1(\register_file.write_data[10] ),
    .A2(_0497_),
    .B1(_0499_),
    .B2(debug_reg3[10]),
    .X(_0119_));
 sky130_fd_sc_hd__a22o_2 _1506_ (.A1(\register_file.write_data[11] ),
    .A2(_0497_),
    .B1(_0499_),
    .B2(debug_reg3[11]),
    .X(_0120_));
 sky130_fd_sc_hd__buf_1 _1507_ (.A(_0496_),
    .X(_0500_));
 sky130_fd_sc_hd__buf_1 _1508_ (.A(_0498_),
    .X(_0501_));
 sky130_fd_sc_hd__a22o_2 _1509_ (.A1(\register_file.write_data[12] ),
    .A2(_0500_),
    .B1(_0501_),
    .B2(debug_reg3[12]),
    .X(_0121_));
 sky130_fd_sc_hd__a22o_2 _1510_ (.A1(\register_file.write_data[13] ),
    .A2(_0500_),
    .B1(_0501_),
    .B2(debug_reg3[13]),
    .X(_0122_));
 sky130_fd_sc_hd__a22o_2 _1511_ (.A1(\register_file.write_data[14] ),
    .A2(_0500_),
    .B1(_0501_),
    .B2(debug_reg3[14]),
    .X(_0123_));
 sky130_fd_sc_hd__a22o_2 _1512_ (.A1(\register_file.write_data[15] ),
    .A2(_0500_),
    .B1(_0501_),
    .B2(debug_reg3[15]),
    .X(_0124_));
 sky130_fd_sc_hd__a22o_2 _1513_ (.A1(\register_file.write_data[16] ),
    .A2(_0500_),
    .B1(_0501_),
    .B2(debug_reg3[16]),
    .X(_0125_));
 sky130_fd_sc_hd__a22o_2 _1514_ (.A1(\register_file.write_data[17] ),
    .A2(_0500_),
    .B1(_0501_),
    .B2(debug_reg3[17]),
    .X(_0126_));
 sky130_fd_sc_hd__a22o_2 _1515_ (.A1(\register_file.write_data[18] ),
    .A2(_0500_),
    .B1(_0501_),
    .B2(debug_reg3[18]),
    .X(_0127_));
 sky130_fd_sc_hd__a22o_2 _1516_ (.A1(\register_file.write_data[19] ),
    .A2(_0500_),
    .B1(_0501_),
    .B2(debug_reg3[19]),
    .X(_0128_));
 sky130_fd_sc_hd__a22o_2 _1517_ (.A1(\register_file.write_data[20] ),
    .A2(_0500_),
    .B1(_0501_),
    .B2(debug_reg3[20]),
    .X(_0129_));
 sky130_fd_sc_hd__a22o_2 _1518_ (.A1(\register_file.write_data[21] ),
    .A2(_0500_),
    .B1(_0501_),
    .B2(debug_reg3[21]),
    .X(_0130_));
 sky130_fd_sc_hd__a22o_2 _1519_ (.A1(\register_file.write_data[22] ),
    .A2(_0500_),
    .B1(_0501_),
    .B2(debug_reg3[22]),
    .X(_0131_));
 sky130_fd_sc_hd__a22o_2 _1520_ (.A1(\register_file.write_data[23] ),
    .A2(_0500_),
    .B1(_0501_),
    .B2(debug_reg3[23]),
    .X(_0132_));
 sky130_fd_sc_hd__a22o_2 _1521_ (.A1(\register_file.write_data[24] ),
    .A2(_0496_),
    .B1(_0498_),
    .B2(debug_reg3[24]),
    .X(_0133_));
 sky130_fd_sc_hd__a22o_2 _1522_ (.A1(\register_file.write_data[25] ),
    .A2(_0496_),
    .B1(_0498_),
    .B2(debug_reg3[25]),
    .X(_0134_));
 sky130_fd_sc_hd__a22o_2 _1523_ (.A1(\register_file.write_data[26] ),
    .A2(_0496_),
    .B1(_0498_),
    .B2(debug_reg3[26]),
    .X(_0135_));
 sky130_fd_sc_hd__a22o_2 _1524_ (.A1(\register_file.write_data[27] ),
    .A2(_0496_),
    .B1(_0498_),
    .B2(debug_reg3[27]),
    .X(_0136_));
 sky130_fd_sc_hd__a22o_2 _1525_ (.A1(\register_file.write_data[28] ),
    .A2(_0496_),
    .B1(_0498_),
    .B2(debug_reg3[28]),
    .X(_0137_));
 sky130_fd_sc_hd__a22o_2 _1526_ (.A1(\register_file.write_data[29] ),
    .A2(_0496_),
    .B1(_0498_),
    .B2(debug_reg3[29]),
    .X(_0138_));
 sky130_fd_sc_hd__a22o_2 _1527_ (.A1(\register_file.write_data[30] ),
    .A2(_0496_),
    .B1(_0498_),
    .B2(debug_reg3[30]),
    .X(_0139_));
 sky130_fd_sc_hd__a22o_2 _1528_ (.A1(\register_file.write_data[31] ),
    .A2(_0496_),
    .B1(_0498_),
    .B2(debug_reg3[31]),
    .X(_0140_));
 sky130_fd_sc_hd__nor3b_2 _1529_ (.A(instruction_debug[22]),
    .B(instruction_debug[23]),
    .C_N(_0071_),
    .Y(_0502_));
 sky130_fd_sc_hd__buf_1 _1530_ (.A(_0502_),
    .X(_0503_));
 sky130_fd_sc_hd__and2_2 _1531_ (.A(debug_reg2[0]),
    .B(_0503_),
    .X(_0141_));
 sky130_fd_sc_hd__and2_2 _1532_ (.A(debug_reg2[1]),
    .B(_0503_),
    .X(_0142_));
 sky130_fd_sc_hd__and2_2 _1533_ (.A(debug_reg2[2]),
    .B(_0503_),
    .X(_0143_));
 sky130_fd_sc_hd__and2_2 _1534_ (.A(debug_reg2[3]),
    .B(_0503_),
    .X(_0144_));
 sky130_fd_sc_hd__and2_2 _1535_ (.A(debug_reg2[4]),
    .B(_0503_),
    .X(_0145_));
 sky130_fd_sc_hd__and2_2 _1536_ (.A(debug_reg2[5]),
    .B(_0503_),
    .X(_0146_));
 sky130_fd_sc_hd__and2_2 _1537_ (.A(debug_reg2[6]),
    .B(_0503_),
    .X(_0147_));
 sky130_fd_sc_hd__and2_2 _1538_ (.A(debug_reg2[7]),
    .B(_0503_),
    .X(_0148_));
 sky130_fd_sc_hd__and2_2 _1539_ (.A(debug_reg2[8]),
    .B(_0503_),
    .X(_0149_));
 sky130_fd_sc_hd__and2_2 _1540_ (.A(debug_reg2[9]),
    .B(_0503_),
    .X(_0150_));
 sky130_fd_sc_hd__and2_2 _1541_ (.A(debug_reg2[10]),
    .B(_0503_),
    .X(_0151_));
 sky130_fd_sc_hd__and2_2 _1542_ (.A(debug_reg2[11]),
    .B(_0503_),
    .X(_0152_));
 sky130_fd_sc_hd__buf_1 _1543_ (.A(_0502_),
    .X(_0504_));
 sky130_fd_sc_hd__and2_2 _1544_ (.A(debug_reg2[12]),
    .B(_0504_),
    .X(_0153_));
 sky130_fd_sc_hd__and2_2 _1545_ (.A(debug_reg2[13]),
    .B(_0504_),
    .X(_0154_));
 sky130_fd_sc_hd__and2_2 _1546_ (.A(debug_reg2[14]),
    .B(_0504_),
    .X(_0155_));
 sky130_fd_sc_hd__and2_2 _1547_ (.A(debug_reg2[15]),
    .B(_0504_),
    .X(_0156_));
 sky130_fd_sc_hd__and2_2 _1548_ (.A(debug_reg2[16]),
    .B(_0504_),
    .X(_0157_));
 sky130_fd_sc_hd__and2_2 _1549_ (.A(debug_reg2[17]),
    .B(_0504_),
    .X(_0158_));
 sky130_fd_sc_hd__and2_2 _1550_ (.A(debug_reg2[18]),
    .B(_0504_),
    .X(_0159_));
 sky130_fd_sc_hd__and2_2 _1551_ (.A(debug_reg2[19]),
    .B(_0504_),
    .X(_0160_));
 sky130_fd_sc_hd__and2_2 _1552_ (.A(debug_reg2[20]),
    .B(_0504_),
    .X(_0161_));
 sky130_fd_sc_hd__and2_2 _1553_ (.A(debug_reg2[21]),
    .B(_0504_),
    .X(_0162_));
 sky130_fd_sc_hd__and2_2 _1554_ (.A(debug_reg2[22]),
    .B(_0504_),
    .X(_0163_));
 sky130_fd_sc_hd__and2_2 _1555_ (.A(debug_reg2[23]),
    .B(_0504_),
    .X(_0164_));
 sky130_fd_sc_hd__and2_2 _1556_ (.A(debug_reg2[24]),
    .B(_0502_),
    .X(_0165_));
 sky130_fd_sc_hd__and2_2 _1557_ (.A(debug_reg2[25]),
    .B(_0502_),
    .X(_0166_));
 sky130_fd_sc_hd__and2_2 _1558_ (.A(debug_reg2[26]),
    .B(_0502_),
    .X(_0167_));
 sky130_fd_sc_hd__and2_2 _1559_ (.A(debug_reg2[27]),
    .B(_0502_),
    .X(_0168_));
 sky130_fd_sc_hd__and2_2 _1560_ (.A(debug_reg2[28]),
    .B(_0502_),
    .X(_0169_));
 sky130_fd_sc_hd__and2_2 _1561_ (.A(debug_reg2[29]),
    .B(_0502_),
    .X(_0170_));
 sky130_fd_sc_hd__and2_2 _1562_ (.A(debug_reg2[30]),
    .B(_0502_),
    .X(_0171_));
 sky130_fd_sc_hd__and2_2 _1563_ (.A(debug_reg2[31]),
    .B(_0502_),
    .X(_0172_));
 sky130_fd_sc_hd__nor2_2 _1564_ (.A(\forwarding_unit.rd_wb[0] ),
    .B(_0493_),
    .Y(_0505_));
 sky130_fd_sc_hd__buf_1 _1565_ (.A(_0505_),
    .X(_0506_));
 sky130_fd_sc_hd__nor2_2 _1566_ (.A(_0521_),
    .B(_0505_),
    .Y(_0507_));
 sky130_fd_sc_hd__buf_1 _1567_ (.A(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__a22o_2 _1568_ (.A1(\register_file.write_data[0] ),
    .A2(_0506_),
    .B1(_0508_),
    .B2(debug_reg2[0]),
    .X(_0173_));
 sky130_fd_sc_hd__a22o_2 _1569_ (.A1(\register_file.write_data[1] ),
    .A2(_0506_),
    .B1(_0508_),
    .B2(debug_reg2[1]),
    .X(_0174_));
 sky130_fd_sc_hd__a22o_2 _1570_ (.A1(\register_file.write_data[2] ),
    .A2(_0506_),
    .B1(_0508_),
    .B2(debug_reg2[2]),
    .X(_0175_));
 sky130_fd_sc_hd__a22o_2 _1571_ (.A1(\register_file.write_data[3] ),
    .A2(_0506_),
    .B1(_0508_),
    .B2(debug_reg2[3]),
    .X(_0176_));
 sky130_fd_sc_hd__a22o_2 _1572_ (.A1(\register_file.write_data[4] ),
    .A2(_0506_),
    .B1(_0508_),
    .B2(debug_reg2[4]),
    .X(_0177_));
 sky130_fd_sc_hd__a22o_2 _1573_ (.A1(\register_file.write_data[5] ),
    .A2(_0506_),
    .B1(_0508_),
    .B2(debug_reg2[5]),
    .X(_0178_));
 sky130_fd_sc_hd__a22o_2 _1574_ (.A1(\register_file.write_data[6] ),
    .A2(_0506_),
    .B1(_0508_),
    .B2(debug_reg2[6]),
    .X(_0179_));
 sky130_fd_sc_hd__a22o_2 _1575_ (.A1(\register_file.write_data[7] ),
    .A2(_0506_),
    .B1(_0508_),
    .B2(debug_reg2[7]),
    .X(_0180_));
 sky130_fd_sc_hd__a22o_2 _1576_ (.A1(\register_file.write_data[8] ),
    .A2(_0506_),
    .B1(_0508_),
    .B2(debug_reg2[8]),
    .X(_0181_));
 sky130_fd_sc_hd__a22o_2 _1577_ (.A1(\register_file.write_data[9] ),
    .A2(_0506_),
    .B1(_0508_),
    .B2(debug_reg2[9]),
    .X(_0182_));
 sky130_fd_sc_hd__a22o_2 _1578_ (.A1(\register_file.write_data[10] ),
    .A2(_0506_),
    .B1(_0508_),
    .B2(debug_reg2[10]),
    .X(_0183_));
 sky130_fd_sc_hd__a22o_2 _1579_ (.A1(\register_file.write_data[11] ),
    .A2(_0506_),
    .B1(_0508_),
    .B2(debug_reg2[11]),
    .X(_0184_));
 sky130_fd_sc_hd__buf_1 _1580_ (.A(_0505_),
    .X(_0509_));
 sky130_fd_sc_hd__buf_1 _1581_ (.A(_0507_),
    .X(_0510_));
 sky130_fd_sc_hd__a22o_2 _1582_ (.A1(\register_file.write_data[12] ),
    .A2(_0509_),
    .B1(_0510_),
    .B2(debug_reg2[12]),
    .X(_0185_));
 sky130_fd_sc_hd__a22o_2 _1583_ (.A1(\register_file.write_data[13] ),
    .A2(_0509_),
    .B1(_0510_),
    .B2(debug_reg2[13]),
    .X(_0186_));
 sky130_fd_sc_hd__a22o_2 _1584_ (.A1(\register_file.write_data[14] ),
    .A2(_0509_),
    .B1(_0510_),
    .B2(debug_reg2[14]),
    .X(_0187_));
 sky130_fd_sc_hd__a22o_2 _1585_ (.A1(\register_file.write_data[15] ),
    .A2(_0509_),
    .B1(_0510_),
    .B2(debug_reg2[15]),
    .X(_0188_));
 sky130_fd_sc_hd__a22o_2 _1586_ (.A1(\register_file.write_data[16] ),
    .A2(_0509_),
    .B1(_0510_),
    .B2(debug_reg2[16]),
    .X(_0189_));
 sky130_fd_sc_hd__a22o_2 _1587_ (.A1(\register_file.write_data[17] ),
    .A2(_0509_),
    .B1(_0510_),
    .B2(debug_reg2[17]),
    .X(_0190_));
 sky130_fd_sc_hd__a22o_2 _1588_ (.A1(\register_file.write_data[18] ),
    .A2(_0509_),
    .B1(_0510_),
    .B2(debug_reg2[18]),
    .X(_0191_));
 sky130_fd_sc_hd__a22o_2 _1589_ (.A1(\register_file.write_data[19] ),
    .A2(_0509_),
    .B1(_0510_),
    .B2(debug_reg2[19]),
    .X(_0192_));
 sky130_fd_sc_hd__a22o_2 _1590_ (.A1(\register_file.write_data[20] ),
    .A2(_0509_),
    .B1(_0510_),
    .B2(debug_reg2[20]),
    .X(_0193_));
 sky130_fd_sc_hd__a22o_2 _1591_ (.A1(\register_file.write_data[21] ),
    .A2(_0509_),
    .B1(_0510_),
    .B2(debug_reg2[21]),
    .X(_0194_));
 sky130_fd_sc_hd__a22o_2 _1592_ (.A1(\register_file.write_data[22] ),
    .A2(_0509_),
    .B1(_0510_),
    .B2(debug_reg2[22]),
    .X(_0195_));
 sky130_fd_sc_hd__a22o_2 _1593_ (.A1(\register_file.write_data[23] ),
    .A2(_0509_),
    .B1(_0510_),
    .B2(debug_reg2[23]),
    .X(_0196_));
 sky130_fd_sc_hd__a22o_2 _1594_ (.A1(\register_file.write_data[24] ),
    .A2(_0505_),
    .B1(_0507_),
    .B2(debug_reg2[24]),
    .X(_0197_));
 sky130_fd_sc_hd__a22o_2 _1595_ (.A1(\register_file.write_data[25] ),
    .A2(_0505_),
    .B1(_0507_),
    .B2(debug_reg2[25]),
    .X(_0198_));
 sky130_fd_sc_hd__a22o_2 _1596_ (.A1(\register_file.write_data[26] ),
    .A2(_0505_),
    .B1(_0507_),
    .B2(debug_reg2[26]),
    .X(_0199_));
 sky130_fd_sc_hd__a22o_2 _1597_ (.A1(\register_file.write_data[27] ),
    .A2(_0505_),
    .B1(_0507_),
    .B2(debug_reg2[27]),
    .X(_0200_));
 sky130_fd_sc_hd__a22o_2 _1598_ (.A1(\register_file.write_data[28] ),
    .A2(_0505_),
    .B1(_0507_),
    .B2(debug_reg2[28]),
    .X(_0201_));
 sky130_fd_sc_hd__a22o_2 _1599_ (.A1(\register_file.write_data[29] ),
    .A2(_0505_),
    .B1(_0507_),
    .B2(debug_reg2[29]),
    .X(_0202_));
 sky130_fd_sc_hd__a22o_2 _1600_ (.A1(\register_file.write_data[30] ),
    .A2(_0505_),
    .B1(_0507_),
    .B2(debug_reg2[30]),
    .X(_0203_));
 sky130_fd_sc_hd__a22o_2 _1601_ (.A1(\register_file.write_data[31] ),
    .A2(_0505_),
    .B1(_0507_),
    .B2(debug_reg2[31]),
    .X(_0204_));
 sky130_fd_sc_hd__nor2_2 _1602_ (.A(\forwarding_unit.rd_wb[1] ),
    .B(_0493_),
    .Y(_0511_));
 sky130_fd_sc_hd__buf_1 _1603_ (.A(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__nor2_2 _1604_ (.A(_0521_),
    .B(_0511_),
    .Y(_0513_));
 sky130_fd_sc_hd__buf_1 _1605_ (.A(_0513_),
    .X(_0514_));
 sky130_fd_sc_hd__a22o_2 _1606_ (.A1(\register_file.write_data[0] ),
    .A2(_0512_),
    .B1(_0514_),
    .B2(debug_reg1[0]),
    .X(_0205_));
 sky130_fd_sc_hd__a22o_2 _1607_ (.A1(\register_file.write_data[1] ),
    .A2(_0512_),
    .B1(_0514_),
    .B2(debug_reg1[1]),
    .X(_0206_));
 sky130_fd_sc_hd__a22o_2 _1608_ (.A1(\register_file.write_data[2] ),
    .A2(_0512_),
    .B1(_0514_),
    .B2(debug_reg1[2]),
    .X(_0207_));
 sky130_fd_sc_hd__a22o_2 _1609_ (.A1(\register_file.write_data[3] ),
    .A2(_0512_),
    .B1(_0514_),
    .B2(debug_reg1[3]),
    .X(_0208_));
 sky130_fd_sc_hd__a22o_2 _1610_ (.A1(\register_file.write_data[4] ),
    .A2(_0512_),
    .B1(_0514_),
    .B2(debug_reg1[4]),
    .X(_0209_));
 sky130_fd_sc_hd__a22o_2 _1611_ (.A1(\register_file.write_data[5] ),
    .A2(_0512_),
    .B1(_0514_),
    .B2(debug_reg1[5]),
    .X(_0210_));
 sky130_fd_sc_hd__a22o_2 _1612_ (.A1(\register_file.write_data[6] ),
    .A2(_0512_),
    .B1(_0514_),
    .B2(debug_reg1[6]),
    .X(_0211_));
 sky130_fd_sc_hd__a22o_2 _1613_ (.A1(\register_file.write_data[7] ),
    .A2(_0512_),
    .B1(_0514_),
    .B2(debug_reg1[7]),
    .X(_0212_));
 sky130_fd_sc_hd__a22o_2 _1614_ (.A1(\register_file.write_data[8] ),
    .A2(_0512_),
    .B1(_0514_),
    .B2(debug_reg1[8]),
    .X(_0213_));
 sky130_fd_sc_hd__a22o_2 _1615_ (.A1(\register_file.write_data[9] ),
    .A2(_0512_),
    .B1(_0514_),
    .B2(debug_reg1[9]),
    .X(_0214_));
 sky130_fd_sc_hd__a22o_2 _1616_ (.A1(\register_file.write_data[10] ),
    .A2(_0512_),
    .B1(_0514_),
    .B2(debug_reg1[10]),
    .X(_0215_));
 sky130_fd_sc_hd__a22o_2 _1617_ (.A1(\register_file.write_data[11] ),
    .A2(_0512_),
    .B1(_0514_),
    .B2(debug_reg1[11]),
    .X(_0216_));
 sky130_fd_sc_hd__buf_1 _1618_ (.A(_0511_),
    .X(_0515_));
 sky130_fd_sc_hd__buf_1 _1619_ (.A(_0513_),
    .X(_0516_));
 sky130_fd_sc_hd__a22o_2 _1620_ (.A1(\register_file.write_data[12] ),
    .A2(_0515_),
    .B1(_0516_),
    .B2(debug_reg1[12]),
    .X(_0217_));
 sky130_fd_sc_hd__a22o_2 _1621_ (.A1(\register_file.write_data[13] ),
    .A2(_0515_),
    .B1(_0516_),
    .B2(debug_reg1[13]),
    .X(_0218_));
 sky130_fd_sc_hd__a22o_2 _1622_ (.A1(\register_file.write_data[14] ),
    .A2(_0515_),
    .B1(_0516_),
    .B2(debug_reg1[14]),
    .X(_0219_));
 sky130_fd_sc_hd__a22o_2 _1623_ (.A1(\register_file.write_data[15] ),
    .A2(_0515_),
    .B1(_0516_),
    .B2(debug_reg1[15]),
    .X(_0220_));
 sky130_fd_sc_hd__a22o_2 _1624_ (.A1(\register_file.write_data[16] ),
    .A2(_0515_),
    .B1(_0516_),
    .B2(debug_reg1[16]),
    .X(_0221_));
 sky130_fd_sc_hd__a22o_2 _1625_ (.A1(\register_file.write_data[17] ),
    .A2(_0515_),
    .B1(_0516_),
    .B2(debug_reg1[17]),
    .X(_0222_));
 sky130_fd_sc_hd__a22o_2 _1626_ (.A1(\register_file.write_data[18] ),
    .A2(_0515_),
    .B1(_0516_),
    .B2(debug_reg1[18]),
    .X(_0223_));
 sky130_fd_sc_hd__a22o_2 _1627_ (.A1(\register_file.write_data[19] ),
    .A2(_0515_),
    .B1(_0516_),
    .B2(debug_reg1[19]),
    .X(_0224_));
 sky130_fd_sc_hd__a22o_2 _1628_ (.A1(\register_file.write_data[20] ),
    .A2(_0515_),
    .B1(_0516_),
    .B2(debug_reg1[20]),
    .X(_0225_));
 sky130_fd_sc_hd__a22o_2 _1629_ (.A1(\register_file.write_data[21] ),
    .A2(_0515_),
    .B1(_0516_),
    .B2(debug_reg1[21]),
    .X(_0226_));
 sky130_fd_sc_hd__a22o_2 _1630_ (.A1(\register_file.write_data[22] ),
    .A2(_0515_),
    .B1(_0516_),
    .B2(debug_reg1[22]),
    .X(_0227_));
 sky130_fd_sc_hd__a22o_2 _1631_ (.A1(\register_file.write_data[23] ),
    .A2(_0515_),
    .B1(_0516_),
    .B2(debug_reg1[23]),
    .X(_0228_));
 sky130_fd_sc_hd__a22o_2 _1632_ (.A1(\register_file.write_data[24] ),
    .A2(_0511_),
    .B1(_0513_),
    .B2(debug_reg1[24]),
    .X(_0229_));
 sky130_fd_sc_hd__a22o_2 _1633_ (.A1(\register_file.write_data[25] ),
    .A2(_0511_),
    .B1(_0513_),
    .B2(debug_reg1[25]),
    .X(_0230_));
 sky130_fd_sc_hd__a22o_2 _1634_ (.A1(\register_file.write_data[26] ),
    .A2(_0511_),
    .B1(_0513_),
    .B2(debug_reg1[26]),
    .X(_0231_));
 sky130_fd_sc_hd__a22o_2 _1635_ (.A1(\register_file.write_data[27] ),
    .A2(_0511_),
    .B1(_0513_),
    .B2(debug_reg1[27]),
    .X(_0232_));
 sky130_fd_sc_hd__a22o_2 _1636_ (.A1(\register_file.write_data[28] ),
    .A2(_0511_),
    .B1(_0513_),
    .B2(debug_reg1[28]),
    .X(_0233_));
 sky130_fd_sc_hd__a22o_2 _1637_ (.A1(\register_file.write_data[29] ),
    .A2(_0511_),
    .B1(_0513_),
    .B2(debug_reg1[29]),
    .X(_0234_));
 sky130_fd_sc_hd__a22o_2 _1638_ (.A1(\register_file.write_data[30] ),
    .A2(_0511_),
    .B1(_0513_),
    .B2(debug_reg1[30]),
    .X(_0235_));
 sky130_fd_sc_hd__a22o_2 _1639_ (.A1(\register_file.write_data[31] ),
    .A2(_0511_),
    .B1(_0513_),
    .B2(debug_reg1[31]),
    .X(_0236_));
 sky130_fd_sc_hd__and2_2 _1640_ (.A(_0442_),
    .B(id_reg_write),
    .X(_0237_));
 sky130_fd_sc_hd__inv_2 _1641_ (.A(_0522_),
    .Y(_0238_));
 sky130_fd_sc_hd__nor2_2 _1642_ (.A(instruction_debug[15]),
    .B(_0521_),
    .Y(_0239_));
 sky130_fd_sc_hd__and3_2 _1643_ (.A(_0441_),
    .B(_0411_),
    .C(debug_reg1[0]),
    .X(_0240_));
 sky130_fd_sc_hd__and3_2 _1644_ (.A(_0441_),
    .B(_0411_),
    .C(debug_reg1[1]),
    .X(_0241_));
 sky130_fd_sc_hd__and3_2 _1645_ (.A(_0441_),
    .B(_0411_),
    .C(debug_reg1[2]),
    .X(_0242_));
 sky130_fd_sc_hd__and3_2 _1646_ (.A(_0441_),
    .B(_0411_),
    .C(debug_reg1[3]),
    .X(_0243_));
 sky130_fd_sc_hd__and3_2 _1647_ (.A(_0441_),
    .B(_0411_),
    .C(debug_reg1[4]),
    .X(_0244_));
 sky130_fd_sc_hd__and3_2 _1648_ (.A(_0441_),
    .B(_0411_),
    .C(debug_reg1[5]),
    .X(_0245_));
 sky130_fd_sc_hd__and3_2 _1649_ (.A(_0441_),
    .B(_0411_),
    .C(debug_reg1[6]),
    .X(_0246_));
 sky130_fd_sc_hd__and3_2 _1650_ (.A(_0441_),
    .B(_0411_),
    .C(debug_reg1[7]),
    .X(_0247_));
 sky130_fd_sc_hd__and3_2 _1651_ (.A(_0441_),
    .B(_0411_),
    .C(debug_reg1[8]),
    .X(_0248_));
 sky130_fd_sc_hd__and3_2 _1652_ (.A(_0441_),
    .B(_0411_),
    .C(debug_reg1[9]),
    .X(_0249_));
 sky130_fd_sc_hd__and3_2 _1653_ (.A(_0441_),
    .B(_0411_),
    .C(debug_reg1[10]),
    .X(_0250_));
 sky130_fd_sc_hd__buf_1 _1654_ (.A(instruction_debug[15]),
    .X(_0517_));
 sky130_fd_sc_hd__buf_1 _1655_ (.A(_0519_),
    .X(_0518_));
 sky130_fd_sc_hd__and3_2 _1656_ (.A(_0517_),
    .B(_0518_),
    .C(debug_reg1[11]),
    .X(_0251_));
 sky130_fd_sc_hd__and3_2 _1657_ (.A(_0517_),
    .B(_0518_),
    .C(debug_reg1[12]),
    .X(_0252_));
 sky130_fd_sc_hd__and3_2 _1658_ (.A(_0517_),
    .B(_0518_),
    .C(debug_reg1[13]),
    .X(_0253_));
 sky130_fd_sc_hd__and3_2 _1659_ (.A(_0517_),
    .B(_0518_),
    .C(debug_reg1[14]),
    .X(_0254_));
 sky130_fd_sc_hd__and3_2 _1660_ (.A(_0517_),
    .B(_0518_),
    .C(debug_reg1[15]),
    .X(_0255_));
 sky130_fd_sc_hd__and3_2 _1661_ (.A(_0517_),
    .B(_0518_),
    .C(debug_reg1[16]),
    .X(_0256_));
 sky130_fd_sc_hd__and3_2 _1662_ (.A(_0517_),
    .B(_0518_),
    .C(debug_reg1[17]),
    .X(_0257_));
 sky130_fd_sc_hd__and3_2 _1663_ (.A(_0517_),
    .B(_0518_),
    .C(debug_reg1[18]),
    .X(_0258_));
 sky130_fd_sc_hd__and3_2 _1664_ (.A(_0517_),
    .B(_0518_),
    .C(debug_reg1[19]),
    .X(_0259_));
 sky130_fd_sc_hd__and3_2 _1665_ (.A(_0517_),
    .B(_0518_),
    .C(debug_reg1[20]),
    .X(_0260_));
 sky130_fd_sc_hd__and3_2 _1666_ (.A(_0517_),
    .B(_0518_),
    .C(debug_reg1[21]),
    .X(_0261_));
 sky130_fd_sc_hd__and3_2 _1667_ (.A(_0517_),
    .B(_0518_),
    .C(debug_reg1[22]),
    .X(_0262_));
 sky130_fd_sc_hd__and3_2 _1668_ (.A(instruction_debug[15]),
    .B(_0592_),
    .C(debug_reg1[23]),
    .X(_0263_));
 sky130_fd_sc_hd__and3_2 _1669_ (.A(instruction_debug[15]),
    .B(_0592_),
    .C(debug_reg1[24]),
    .X(_0264_));
 sky130_fd_sc_hd__and3_2 _1670_ (.A(instruction_debug[15]),
    .B(_0592_),
    .C(debug_reg1[25]),
    .X(_0265_));
 sky130_fd_sc_hd__and3_2 _1671_ (.A(instruction_debug[15]),
    .B(_0592_),
    .C(debug_reg1[26]),
    .X(_0266_));
 sky130_fd_sc_hd__and3_2 _1672_ (.A(instruction_debug[15]),
    .B(_0592_),
    .C(debug_reg1[27]),
    .X(_0267_));
 sky130_fd_sc_hd__and3_2 _1673_ (.A(instruction_debug[15]),
    .B(_0592_),
    .C(debug_reg1[28]),
    .X(_0268_));
 sky130_fd_sc_hd__and3_2 _1674_ (.A(instruction_debug[15]),
    .B(_0592_),
    .C(debug_reg1[29]),
    .X(_0269_));
 sky130_fd_sc_hd__and3_2 _1675_ (.A(instruction_debug[15]),
    .B(_0592_),
    .C(debug_reg1[30]),
    .X(_0270_));
 sky130_fd_sc_hd__and3_2 _1676_ (.A(instruction_debug[15]),
    .B(_0592_),
    .C(debug_reg1[31]),
    .X(_0271_));
 sky130_fd_sc_hd__and2_2 _1677_ (.A(instruction_debug[21]),
    .B(_0239_),
    .X(_0272_));
 sky130_fd_sc_hd__and2_2 _1678_ (.A(instruction_debug[22]),
    .B(_0239_),
    .X(_0273_));
 sky130_fd_sc_hd__and2_2 _1679_ (.A(instruction_debug[23]),
    .B(_0239_),
    .X(_0274_));
 sky130_fd_sc_hd__nor2_2 _1680_ (.A(pc_current[2]),
    .B(_0440_),
    .Y(_0275_));
 sky130_fd_sc_hd__nor2b_2 _1681_ (.A(_0443_),
    .B_N(_0275_),
    .Y(_0276_));
 sky130_fd_sc_hd__nor2b_2 _1682_ (.A(pc_current[3]),
    .B_N(_0275_),
    .Y(_0277_));
 sky130_fd_sc_hd__nor2_2 _1683_ (.A(_0440_),
    .B(_0443_),
    .Y(_0278_));
 sky130_fd_sc_hd__dfxtp_2 _1684_ (.CLK(clk),
    .D(_0001_),
    .Q(\register_file.write_data[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1685_ (.CLK(clk),
    .D(_0002_),
    .Q(\register_file.write_data[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1686_ (.CLK(clk),
    .D(_0003_),
    .Q(\register_file.write_data[2] ));
 sky130_fd_sc_hd__dfxtp_2 _1687_ (.CLK(clk),
    .D(_0004_),
    .Q(\register_file.write_data[3] ));
 sky130_fd_sc_hd__dfxtp_2 _1688_ (.CLK(clk),
    .D(_0005_),
    .Q(\register_file.write_data[4] ));
 sky130_fd_sc_hd__dfxtp_2 _1689_ (.CLK(clk),
    .D(_0006_),
    .Q(\register_file.write_data[5] ));
 sky130_fd_sc_hd__dfxtp_2 _1690_ (.CLK(clk),
    .D(_0007_),
    .Q(\register_file.write_data[6] ));
 sky130_fd_sc_hd__dfxtp_2 _1691_ (.CLK(clk),
    .D(_0008_),
    .Q(\register_file.write_data[7] ));
 sky130_fd_sc_hd__dfxtp_2 _1692_ (.CLK(clk),
    .D(_0009_),
    .Q(\register_file.write_data[8] ));
 sky130_fd_sc_hd__dfxtp_2 _1693_ (.CLK(clk),
    .D(_0010_),
    .Q(\register_file.write_data[9] ));
 sky130_fd_sc_hd__dfxtp_2 _1694_ (.CLK(clk),
    .D(_0011_),
    .Q(\register_file.write_data[10] ));
 sky130_fd_sc_hd__dfxtp_2 _1695_ (.CLK(clk),
    .D(_0012_),
    .Q(\register_file.write_data[11] ));
 sky130_fd_sc_hd__dfxtp_2 _1696_ (.CLK(clk),
    .D(_0013_),
    .Q(\register_file.write_data[12] ));
 sky130_fd_sc_hd__dfxtp_2 _1697_ (.CLK(clk),
    .D(_0014_),
    .Q(\register_file.write_data[13] ));
 sky130_fd_sc_hd__dfxtp_2 _1698_ (.CLK(clk),
    .D(_0015_),
    .Q(\register_file.write_data[14] ));
 sky130_fd_sc_hd__dfxtp_2 _1699_ (.CLK(clk),
    .D(_0016_),
    .Q(\register_file.write_data[15] ));
 sky130_fd_sc_hd__dfxtp_2 _1700_ (.CLK(clk),
    .D(_0017_),
    .Q(\register_file.write_data[16] ));
 sky130_fd_sc_hd__dfxtp_2 _1701_ (.CLK(clk),
    .D(_0018_),
    .Q(\register_file.write_data[17] ));
 sky130_fd_sc_hd__dfxtp_2 _1702_ (.CLK(clk),
    .D(_0019_),
    .Q(\register_file.write_data[18] ));
 sky130_fd_sc_hd__dfxtp_2 _1703_ (.CLK(clk),
    .D(_0020_),
    .Q(\register_file.write_data[19] ));
 sky130_fd_sc_hd__dfxtp_2 _1704_ (.CLK(clk),
    .D(_0021_),
    .Q(\register_file.write_data[20] ));
 sky130_fd_sc_hd__dfxtp_2 _1705_ (.CLK(clk),
    .D(_0022_),
    .Q(\register_file.write_data[21] ));
 sky130_fd_sc_hd__dfxtp_2 _1706_ (.CLK(clk),
    .D(_0023_),
    .Q(\register_file.write_data[22] ));
 sky130_fd_sc_hd__dfxtp_2 _1707_ (.CLK(clk),
    .D(_0024_),
    .Q(\register_file.write_data[23] ));
 sky130_fd_sc_hd__dfxtp_2 _1708_ (.CLK(clk),
    .D(_0025_),
    .Q(\register_file.write_data[24] ));
 sky130_fd_sc_hd__dfxtp_2 _1709_ (.CLK(clk),
    .D(_0026_),
    .Q(\register_file.write_data[25] ));
 sky130_fd_sc_hd__dfxtp_2 _1710_ (.CLK(clk),
    .D(_0027_),
    .Q(\register_file.write_data[26] ));
 sky130_fd_sc_hd__dfxtp_2 _1711_ (.CLK(clk),
    .D(_0028_),
    .Q(\register_file.write_data[27] ));
 sky130_fd_sc_hd__dfxtp_2 _1712_ (.CLK(clk),
    .D(_0029_),
    .Q(\register_file.write_data[28] ));
 sky130_fd_sc_hd__dfxtp_2 _1713_ (.CLK(clk),
    .D(_0030_),
    .Q(\register_file.write_data[29] ));
 sky130_fd_sc_hd__dfxtp_2 _1714_ (.CLK(clk),
    .D(_0031_),
    .Q(\register_file.write_data[30] ));
 sky130_fd_sc_hd__dfxtp_2 _1715_ (.CLK(clk),
    .D(_0032_),
    .Q(\register_file.write_data[31] ));
 sky130_fd_sc_hd__dfxtp_2 _1716_ (.CLK(clk),
    .D(_0033_),
    .Q(\ex_mem_alu_result[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1717_ (.CLK(clk),
    .D(_0034_),
    .Q(\ex_mem_alu_result[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1718_ (.CLK(clk),
    .D(_0035_),
    .Q(\dmem.address[2] ));
 sky130_fd_sc_hd__dfxtp_2 _1719_ (.CLK(clk),
    .D(_0036_),
    .Q(\dmem.address[3] ));
 sky130_fd_sc_hd__dfxtp_2 _1720_ (.CLK(clk),
    .D(_0037_),
    .Q(\dmem.address[4] ));
 sky130_fd_sc_hd__dfxtp_2 _1721_ (.CLK(clk),
    .D(_0038_),
    .Q(\dmem.address[5] ));
 sky130_fd_sc_hd__dfxtp_2 _1722_ (.CLK(clk),
    .D(_0039_),
    .Q(\dmem.address[6] ));
 sky130_fd_sc_hd__dfxtp_2 _1723_ (.CLK(clk),
    .D(_0040_),
    .Q(\dmem.address[7] ));
 sky130_fd_sc_hd__dfxtp_2 _1724_ (.CLK(clk),
    .D(_0041_),
    .Q(\dmem.address[8] ));
 sky130_fd_sc_hd__dfxtp_2 _1725_ (.CLK(clk),
    .D(_0042_),
    .Q(\dmem.address[9] ));
 sky130_fd_sc_hd__dfxtp_2 _1726_ (.CLK(clk),
    .D(_0043_),
    .Q(\dmem.address[10] ));
 sky130_fd_sc_hd__dfxtp_2 _1727_ (.CLK(clk),
    .D(_0044_),
    .Q(\dmem.address[11] ));
 sky130_fd_sc_hd__dfxtp_2 _1728_ (.CLK(clk),
    .D(_0045_),
    .Q(\dmem.address[12] ));
 sky130_fd_sc_hd__dfxtp_2 _1729_ (.CLK(clk),
    .D(_0046_),
    .Q(\dmem.address[13] ));
 sky130_fd_sc_hd__dfxtp_2 _1730_ (.CLK(clk),
    .D(_0047_),
    .Q(\dmem.address[14] ));
 sky130_fd_sc_hd__dfxtp_2 _1731_ (.CLK(clk),
    .D(_0048_),
    .Q(\dmem.address[15] ));
 sky130_fd_sc_hd__dfxtp_2 _1732_ (.CLK(clk),
    .D(_0049_),
    .Q(\dmem.address[16] ));
 sky130_fd_sc_hd__dfxtp_2 _1733_ (.CLK(clk),
    .D(_0050_),
    .Q(\dmem.address[17] ));
 sky130_fd_sc_hd__dfxtp_2 _1734_ (.CLK(clk),
    .D(_0051_),
    .Q(\dmem.address[18] ));
 sky130_fd_sc_hd__dfxtp_2 _1735_ (.CLK(clk),
    .D(_0052_),
    .Q(\dmem.address[19] ));
 sky130_fd_sc_hd__dfxtp_2 _1736_ (.CLK(clk),
    .D(_0053_),
    .Q(\dmem.address[20] ));
 sky130_fd_sc_hd__dfxtp_2 _1737_ (.CLK(clk),
    .D(_0054_),
    .Q(\dmem.address[21] ));
 sky130_fd_sc_hd__dfxtp_2 _1738_ (.CLK(clk),
    .D(_0055_),
    .Q(\dmem.address[22] ));
 sky130_fd_sc_hd__dfxtp_2 _1739_ (.CLK(clk),
    .D(_0056_),
    .Q(\dmem.address[23] ));
 sky130_fd_sc_hd__dfxtp_2 _1740_ (.CLK(clk),
    .D(_0057_),
    .Q(\dmem.address[24] ));
 sky130_fd_sc_hd__dfxtp_2 _1741_ (.CLK(clk),
    .D(_0058_),
    .Q(\dmem.address[25] ));
 sky130_fd_sc_hd__dfxtp_2 _1742_ (.CLK(clk),
    .D(_0059_),
    .Q(\dmem.address[26] ));
 sky130_fd_sc_hd__dfxtp_2 _1743_ (.CLK(clk),
    .D(_0060_),
    .Q(\dmem.address[27] ));
 sky130_fd_sc_hd__dfxtp_2 _1744_ (.CLK(clk),
    .D(_0061_),
    .Q(\dmem.address[28] ));
 sky130_fd_sc_hd__dfxtp_2 _1745_ (.CLK(clk),
    .D(_0062_),
    .Q(\dmem.address[29] ));
 sky130_fd_sc_hd__dfxtp_2 _1746_ (.CLK(clk),
    .D(_0063_),
    .Q(\dmem.address[30] ));
 sky130_fd_sc_hd__dfxtp_2 _1747_ (.CLK(clk),
    .D(_0064_),
    .Q(\dmem.address[31] ));
 sky130_fd_sc_hd__dfxtp_2 _1748_ (.CLK(clk),
    .D(_0065_),
    .Q(mem_wb_valid));
 sky130_fd_sc_hd__dfxtp_2 _1749_ (.CLK(clk),
    .D(_0066_),
    .Q(ex_mem_valid));
 sky130_fd_sc_hd__dfxtp_2 _1750_ (.CLK(clk),
    .D(_0067_),
    .Q(\forwarding_unit.rd_wb[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1751_ (.CLK(clk),
    .D(_0068_),
    .Q(\forwarding_unit.rd_wb[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1752_ (.CLK(clk),
    .D(_0069_),
    .Q(instruction_debug[23]));
 sky130_fd_sc_hd__dfxtp_2 _1753_ (.CLK(clk),
    .D(_0070_),
    .Q(\forwarding_unit.rs1_ex[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1754_ (.CLK(clk),
    .D(_0071_),
    .Q(\forwarding_unit.rs2_ex[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1755_ (.CLK(clk),
    .D(_0072_),
    .Q(\forwarding_unit.rs2_ex[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1756_ (.CLK(clk),
    .D(_0073_),
    .Q(\forwarding_unit.rs2_ex[3] ));
 sky130_fd_sc_hd__dfxtp_2 _1757_ (.CLK(clk),
    .D(_0074_),
    .Q(\id_ex_rd_addr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1758_ (.CLK(clk),
    .D(_0075_),
    .Q(id_ex_valid));
 sky130_fd_sc_hd__dfxtp_2 _1759_ (.CLK(clk),
    .D(_0000_),
    .Q(if_id_valid));
 sky130_fd_sc_hd__dfxtp_2 _1760_ (.CLK(clk),
    .D(_0076_),
    .Q(\forwarding_unit.rd_mem[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1761_ (.CLK(clk),
    .D(_0077_),
    .Q(\forwarding_unit.rd_mem[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1762_ (.CLK(clk),
    .D(_0078_),
    .Q(\forwarding_unit.reg_write_wb ));
 sky130_fd_sc_hd__dfxtp_2 _1763_ (.CLK(clk),
    .D(_0079_),
    .Q(pc_current[2]));
 sky130_fd_sc_hd__dfxtp_2 _1764_ (.CLK(clk),
    .D(_0080_),
    .Q(pc_current[3]));
 sky130_fd_sc_hd__dfxtp_2 _1765_ (.CLK(clk),
    .D(_0081_),
    .Q(pc_current[4]));
 sky130_fd_sc_hd__dfxtp_2 _1766_ (.CLK(clk),
    .D(_0082_),
    .Q(pc_current[5]));
 sky130_fd_sc_hd__dfxtp_2 _1767_ (.CLK(clk),
    .D(_0083_),
    .Q(pc_current[6]));
 sky130_fd_sc_hd__dfxtp_2 _1768_ (.CLK(clk),
    .D(_0084_),
    .Q(pc_current[7]));
 sky130_fd_sc_hd__dfxtp_2 _1769_ (.CLK(clk),
    .D(_0085_),
    .Q(pc_current[8]));
 sky130_fd_sc_hd__dfxtp_2 _1770_ (.CLK(clk),
    .D(_0086_),
    .Q(pc_current[9]));
 sky130_fd_sc_hd__dfxtp_2 _1771_ (.CLK(clk),
    .D(_0087_),
    .Q(pc_current[10]));
 sky130_fd_sc_hd__dfxtp_2 _1772_ (.CLK(clk),
    .D(_0088_),
    .Q(pc_current[11]));
 sky130_fd_sc_hd__dfxtp_2 _1773_ (.CLK(clk),
    .D(_0089_),
    .Q(pc_current[12]));
 sky130_fd_sc_hd__dfxtp_2 _1774_ (.CLK(clk),
    .D(_0090_),
    .Q(pc_current[13]));
 sky130_fd_sc_hd__dfxtp_2 _1775_ (.CLK(clk),
    .D(_0091_),
    .Q(pc_current[14]));
 sky130_fd_sc_hd__dfxtp_2 _1776_ (.CLK(clk),
    .D(_0092_),
    .Q(pc_current[15]));
 sky130_fd_sc_hd__dfxtp_2 _1777_ (.CLK(clk),
    .D(_0093_),
    .Q(pc_current[16]));
 sky130_fd_sc_hd__dfxtp_2 _1778_ (.CLK(clk),
    .D(_0094_),
    .Q(pc_current[17]));
 sky130_fd_sc_hd__dfxtp_2 _1779_ (.CLK(clk),
    .D(_0095_),
    .Q(pc_current[18]));
 sky130_fd_sc_hd__dfxtp_2 _1780_ (.CLK(clk),
    .D(_0096_),
    .Q(pc_current[19]));
 sky130_fd_sc_hd__dfxtp_2 _1781_ (.CLK(clk),
    .D(_0097_),
    .Q(pc_current[20]));
 sky130_fd_sc_hd__dfxtp_2 _1782_ (.CLK(clk),
    .D(_0098_),
    .Q(pc_current[21]));
 sky130_fd_sc_hd__dfxtp_2 _1783_ (.CLK(clk),
    .D(_0099_),
    .Q(pc_current[22]));
 sky130_fd_sc_hd__dfxtp_2 _1784_ (.CLK(clk),
    .D(_0100_),
    .Q(pc_current[23]));
 sky130_fd_sc_hd__dfxtp_2 _1785_ (.CLK(clk),
    .D(_0101_),
    .Q(pc_current[24]));
 sky130_fd_sc_hd__dfxtp_2 _1786_ (.CLK(clk),
    .D(_0102_),
    .Q(pc_current[25]));
 sky130_fd_sc_hd__dfxtp_2 _1787_ (.CLK(clk),
    .D(_0103_),
    .Q(pc_current[26]));
 sky130_fd_sc_hd__dfxtp_2 _1788_ (.CLK(clk),
    .D(_0104_),
    .Q(pc_current[27]));
 sky130_fd_sc_hd__dfxtp_2 _1789_ (.CLK(clk),
    .D(_0105_),
    .Q(pc_current[28]));
 sky130_fd_sc_hd__dfxtp_2 _1790_ (.CLK(clk),
    .D(_0106_),
    .Q(pc_current[29]));
 sky130_fd_sc_hd__dfxtp_2 _1791_ (.CLK(clk),
    .D(_0107_),
    .Q(pc_current[30]));
 sky130_fd_sc_hd__dfxtp_2 _1792_ (.CLK(clk),
    .D(_0108_),
    .Q(pc_current[31]));
 sky130_fd_sc_hd__dfxtp_2 _1793_ (.CLK(clk),
    .D(_0109_),
    .Q(debug_reg3[0]));
 sky130_fd_sc_hd__dfxtp_2 _1794_ (.CLK(clk),
    .D(_0110_),
    .Q(debug_reg3[1]));
 sky130_fd_sc_hd__dfxtp_2 _1795_ (.CLK(clk),
    .D(_0111_),
    .Q(debug_reg3[2]));
 sky130_fd_sc_hd__dfxtp_2 _1796_ (.CLK(clk),
    .D(_0112_),
    .Q(debug_reg3[3]));
 sky130_fd_sc_hd__dfxtp_2 _1797_ (.CLK(clk),
    .D(_0113_),
    .Q(debug_reg3[4]));
 sky130_fd_sc_hd__dfxtp_2 _1798_ (.CLK(clk),
    .D(_0114_),
    .Q(debug_reg3[5]));
 sky130_fd_sc_hd__dfxtp_2 _1799_ (.CLK(clk),
    .D(_0115_),
    .Q(debug_reg3[6]));
 sky130_fd_sc_hd__dfxtp_2 _1800_ (.CLK(clk),
    .D(_0116_),
    .Q(debug_reg3[7]));
 sky130_fd_sc_hd__dfxtp_2 _1801_ (.CLK(clk),
    .D(_0117_),
    .Q(debug_reg3[8]));
 sky130_fd_sc_hd__dfxtp_2 _1802_ (.CLK(clk),
    .D(_0118_),
    .Q(debug_reg3[9]));
 sky130_fd_sc_hd__dfxtp_2 _1803_ (.CLK(clk),
    .D(_0119_),
    .Q(debug_reg3[10]));
 sky130_fd_sc_hd__dfxtp_2 _1804_ (.CLK(clk),
    .D(_0120_),
    .Q(debug_reg3[11]));
 sky130_fd_sc_hd__dfxtp_2 _1805_ (.CLK(clk),
    .D(_0121_),
    .Q(debug_reg3[12]));
 sky130_fd_sc_hd__dfxtp_2 _1806_ (.CLK(clk),
    .D(_0122_),
    .Q(debug_reg3[13]));
 sky130_fd_sc_hd__dfxtp_2 _1807_ (.CLK(clk),
    .D(_0123_),
    .Q(debug_reg3[14]));
 sky130_fd_sc_hd__dfxtp_2 _1808_ (.CLK(clk),
    .D(_0124_),
    .Q(debug_reg3[15]));
 sky130_fd_sc_hd__dfxtp_2 _1809_ (.CLK(clk),
    .D(_0125_),
    .Q(debug_reg3[16]));
 sky130_fd_sc_hd__dfxtp_2 _1810_ (.CLK(clk),
    .D(_0126_),
    .Q(debug_reg3[17]));
 sky130_fd_sc_hd__dfxtp_2 _1811_ (.CLK(clk),
    .D(_0127_),
    .Q(debug_reg3[18]));
 sky130_fd_sc_hd__dfxtp_2 _1812_ (.CLK(clk),
    .D(_0128_),
    .Q(debug_reg3[19]));
 sky130_fd_sc_hd__dfxtp_2 _1813_ (.CLK(clk),
    .D(_0129_),
    .Q(debug_reg3[20]));
 sky130_fd_sc_hd__dfxtp_2 _1814_ (.CLK(clk),
    .D(_0130_),
    .Q(debug_reg3[21]));
 sky130_fd_sc_hd__dfxtp_2 _1815_ (.CLK(clk),
    .D(_0131_),
    .Q(debug_reg3[22]));
 sky130_fd_sc_hd__dfxtp_2 _1816_ (.CLK(clk),
    .D(_0132_),
    .Q(debug_reg3[23]));
 sky130_fd_sc_hd__dfxtp_2 _1817_ (.CLK(clk),
    .D(_0133_),
    .Q(debug_reg3[24]));
 sky130_fd_sc_hd__dfxtp_2 _1818_ (.CLK(clk),
    .D(_0134_),
    .Q(debug_reg3[25]));
 sky130_fd_sc_hd__dfxtp_2 _1819_ (.CLK(clk),
    .D(_0135_),
    .Q(debug_reg3[26]));
 sky130_fd_sc_hd__dfxtp_2 _1820_ (.CLK(clk),
    .D(_0136_),
    .Q(debug_reg3[27]));
 sky130_fd_sc_hd__dfxtp_2 _1821_ (.CLK(clk),
    .D(_0137_),
    .Q(debug_reg3[28]));
 sky130_fd_sc_hd__dfxtp_2 _1822_ (.CLK(clk),
    .D(_0138_),
    .Q(debug_reg3[29]));
 sky130_fd_sc_hd__dfxtp_2 _1823_ (.CLK(clk),
    .D(_0139_),
    .Q(debug_reg3[30]));
 sky130_fd_sc_hd__dfxtp_2 _1824_ (.CLK(clk),
    .D(_0140_),
    .Q(debug_reg3[31]));
 sky130_fd_sc_hd__dfxtp_2 _1825_ (.CLK(clk),
    .D(_0141_),
    .Q(\id_ex_rs2_data[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1826_ (.CLK(clk),
    .D(_0142_),
    .Q(\id_ex_rs2_data[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1827_ (.CLK(clk),
    .D(_0143_),
    .Q(\id_ex_rs2_data[2] ));
 sky130_fd_sc_hd__dfxtp_2 _1828_ (.CLK(clk),
    .D(_0144_),
    .Q(\id_ex_rs2_data[3] ));
 sky130_fd_sc_hd__dfxtp_2 _1829_ (.CLK(clk),
    .D(_0145_),
    .Q(\id_ex_rs2_data[4] ));
 sky130_fd_sc_hd__dfxtp_2 _1830_ (.CLK(clk),
    .D(_0146_),
    .Q(\id_ex_rs2_data[5] ));
 sky130_fd_sc_hd__dfxtp_2 _1831_ (.CLK(clk),
    .D(_0147_),
    .Q(\id_ex_rs2_data[6] ));
 sky130_fd_sc_hd__dfxtp_2 _1832_ (.CLK(clk),
    .D(_0148_),
    .Q(\id_ex_rs2_data[7] ));
 sky130_fd_sc_hd__dfxtp_2 _1833_ (.CLK(clk),
    .D(_0149_),
    .Q(\id_ex_rs2_data[8] ));
 sky130_fd_sc_hd__dfxtp_2 _1834_ (.CLK(clk),
    .D(_0150_),
    .Q(\id_ex_rs2_data[9] ));
 sky130_fd_sc_hd__dfxtp_2 _1835_ (.CLK(clk),
    .D(_0151_),
    .Q(\id_ex_rs2_data[10] ));
 sky130_fd_sc_hd__dfxtp_2 _1836_ (.CLK(clk),
    .D(_0152_),
    .Q(\id_ex_rs2_data[11] ));
 sky130_fd_sc_hd__dfxtp_2 _1837_ (.CLK(clk),
    .D(_0153_),
    .Q(\id_ex_rs2_data[12] ));
 sky130_fd_sc_hd__dfxtp_2 _1838_ (.CLK(clk),
    .D(_0154_),
    .Q(\id_ex_rs2_data[13] ));
 sky130_fd_sc_hd__dfxtp_2 _1839_ (.CLK(clk),
    .D(_0155_),
    .Q(\id_ex_rs2_data[14] ));
 sky130_fd_sc_hd__dfxtp_2 _1840_ (.CLK(clk),
    .D(_0156_),
    .Q(\id_ex_rs2_data[15] ));
 sky130_fd_sc_hd__dfxtp_2 _1841_ (.CLK(clk),
    .D(_0157_),
    .Q(\id_ex_rs2_data[16] ));
 sky130_fd_sc_hd__dfxtp_2 _1842_ (.CLK(clk),
    .D(_0158_),
    .Q(\id_ex_rs2_data[17] ));
 sky130_fd_sc_hd__dfxtp_2 _1843_ (.CLK(clk),
    .D(_0159_),
    .Q(\id_ex_rs2_data[18] ));
 sky130_fd_sc_hd__dfxtp_2 _1844_ (.CLK(clk),
    .D(_0160_),
    .Q(\id_ex_rs2_data[19] ));
 sky130_fd_sc_hd__dfxtp_2 _1845_ (.CLK(clk),
    .D(_0161_),
    .Q(\id_ex_rs2_data[20] ));
 sky130_fd_sc_hd__dfxtp_2 _1846_ (.CLK(clk),
    .D(_0162_),
    .Q(\id_ex_rs2_data[21] ));
 sky130_fd_sc_hd__dfxtp_2 _1847_ (.CLK(clk),
    .D(_0163_),
    .Q(\id_ex_rs2_data[22] ));
 sky130_fd_sc_hd__dfxtp_2 _1848_ (.CLK(clk),
    .D(_0164_),
    .Q(\id_ex_rs2_data[23] ));
 sky130_fd_sc_hd__dfxtp_2 _1849_ (.CLK(clk),
    .D(_0165_),
    .Q(\id_ex_rs2_data[24] ));
 sky130_fd_sc_hd__dfxtp_2 _1850_ (.CLK(clk),
    .D(_0166_),
    .Q(\id_ex_rs2_data[25] ));
 sky130_fd_sc_hd__dfxtp_2 _1851_ (.CLK(clk),
    .D(_0167_),
    .Q(\id_ex_rs2_data[26] ));
 sky130_fd_sc_hd__dfxtp_2 _1852_ (.CLK(clk),
    .D(_0168_),
    .Q(\id_ex_rs2_data[27] ));
 sky130_fd_sc_hd__dfxtp_2 _1853_ (.CLK(clk),
    .D(_0169_),
    .Q(\id_ex_rs2_data[28] ));
 sky130_fd_sc_hd__dfxtp_2 _1854_ (.CLK(clk),
    .D(_0170_),
    .Q(\id_ex_rs2_data[29] ));
 sky130_fd_sc_hd__dfxtp_2 _1855_ (.CLK(clk),
    .D(_0171_),
    .Q(\id_ex_rs2_data[30] ));
 sky130_fd_sc_hd__dfxtp_2 _1856_ (.CLK(clk),
    .D(_0172_),
    .Q(\id_ex_rs2_data[31] ));
 sky130_fd_sc_hd__dfxtp_2 _1857_ (.CLK(clk),
    .D(_0173_),
    .Q(debug_reg2[0]));
 sky130_fd_sc_hd__dfxtp_2 _1858_ (.CLK(clk),
    .D(_0174_),
    .Q(debug_reg2[1]));
 sky130_fd_sc_hd__dfxtp_2 _1859_ (.CLK(clk),
    .D(_0175_),
    .Q(debug_reg2[2]));
 sky130_fd_sc_hd__dfxtp_2 _1860_ (.CLK(clk),
    .D(_0176_),
    .Q(debug_reg2[3]));
 sky130_fd_sc_hd__dfxtp_2 _1861_ (.CLK(clk),
    .D(_0177_),
    .Q(debug_reg2[4]));
 sky130_fd_sc_hd__dfxtp_2 _1862_ (.CLK(clk),
    .D(_0178_),
    .Q(debug_reg2[5]));
 sky130_fd_sc_hd__dfxtp_2 _1863_ (.CLK(clk),
    .D(_0179_),
    .Q(debug_reg2[6]));
 sky130_fd_sc_hd__dfxtp_2 _1864_ (.CLK(clk),
    .D(_0180_),
    .Q(debug_reg2[7]));
 sky130_fd_sc_hd__dfxtp_2 _1865_ (.CLK(clk),
    .D(_0181_),
    .Q(debug_reg2[8]));
 sky130_fd_sc_hd__dfxtp_2 _1866_ (.CLK(clk),
    .D(_0182_),
    .Q(debug_reg2[9]));
 sky130_fd_sc_hd__dfxtp_2 _1867_ (.CLK(clk),
    .D(_0183_),
    .Q(debug_reg2[10]));
 sky130_fd_sc_hd__dfxtp_2 _1868_ (.CLK(clk),
    .D(_0184_),
    .Q(debug_reg2[11]));
 sky130_fd_sc_hd__dfxtp_2 _1869_ (.CLK(clk),
    .D(_0185_),
    .Q(debug_reg2[12]));
 sky130_fd_sc_hd__dfxtp_2 _1870_ (.CLK(clk),
    .D(_0186_),
    .Q(debug_reg2[13]));
 sky130_fd_sc_hd__dfxtp_2 _1871_ (.CLK(clk),
    .D(_0187_),
    .Q(debug_reg2[14]));
 sky130_fd_sc_hd__dfxtp_2 _1872_ (.CLK(clk),
    .D(_0188_),
    .Q(debug_reg2[15]));
 sky130_fd_sc_hd__dfxtp_2 _1873_ (.CLK(clk),
    .D(_0189_),
    .Q(debug_reg2[16]));
 sky130_fd_sc_hd__dfxtp_2 _1874_ (.CLK(clk),
    .D(_0190_),
    .Q(debug_reg2[17]));
 sky130_fd_sc_hd__dfxtp_2 _1875_ (.CLK(clk),
    .D(_0191_),
    .Q(debug_reg2[18]));
 sky130_fd_sc_hd__dfxtp_2 _1876_ (.CLK(clk),
    .D(_0192_),
    .Q(debug_reg2[19]));
 sky130_fd_sc_hd__dfxtp_2 _1877_ (.CLK(clk),
    .D(_0193_),
    .Q(debug_reg2[20]));
 sky130_fd_sc_hd__dfxtp_2 _1878_ (.CLK(clk),
    .D(_0194_),
    .Q(debug_reg2[21]));
 sky130_fd_sc_hd__dfxtp_2 _1879_ (.CLK(clk),
    .D(_0195_),
    .Q(debug_reg2[22]));
 sky130_fd_sc_hd__dfxtp_2 _1880_ (.CLK(clk),
    .D(_0196_),
    .Q(debug_reg2[23]));
 sky130_fd_sc_hd__dfxtp_2 _1881_ (.CLK(clk),
    .D(_0197_),
    .Q(debug_reg2[24]));
 sky130_fd_sc_hd__dfxtp_2 _1882_ (.CLK(clk),
    .D(_0198_),
    .Q(debug_reg2[25]));
 sky130_fd_sc_hd__dfxtp_2 _1883_ (.CLK(clk),
    .D(_0199_),
    .Q(debug_reg2[26]));
 sky130_fd_sc_hd__dfxtp_2 _1884_ (.CLK(clk),
    .D(_0200_),
    .Q(debug_reg2[27]));
 sky130_fd_sc_hd__dfxtp_2 _1885_ (.CLK(clk),
    .D(_0201_),
    .Q(debug_reg2[28]));
 sky130_fd_sc_hd__dfxtp_2 _1886_ (.CLK(clk),
    .D(_0202_),
    .Q(debug_reg2[29]));
 sky130_fd_sc_hd__dfxtp_2 _1887_ (.CLK(clk),
    .D(_0203_),
    .Q(debug_reg2[30]));
 sky130_fd_sc_hd__dfxtp_2 _1888_ (.CLK(clk),
    .D(_0204_),
    .Q(debug_reg2[31]));
 sky130_fd_sc_hd__dfxtp_2 _1889_ (.CLK(clk),
    .D(_0205_),
    .Q(debug_reg1[0]));
 sky130_fd_sc_hd__dfxtp_2 _1890_ (.CLK(clk),
    .D(_0206_),
    .Q(debug_reg1[1]));
 sky130_fd_sc_hd__dfxtp_2 _1891_ (.CLK(clk),
    .D(_0207_),
    .Q(debug_reg1[2]));
 sky130_fd_sc_hd__dfxtp_2 _1892_ (.CLK(clk),
    .D(_0208_),
    .Q(debug_reg1[3]));
 sky130_fd_sc_hd__dfxtp_2 _1893_ (.CLK(clk),
    .D(_0209_),
    .Q(debug_reg1[4]));
 sky130_fd_sc_hd__dfxtp_2 _1894_ (.CLK(clk),
    .D(_0210_),
    .Q(debug_reg1[5]));
 sky130_fd_sc_hd__dfxtp_2 _1895_ (.CLK(clk),
    .D(_0211_),
    .Q(debug_reg1[6]));
 sky130_fd_sc_hd__dfxtp_2 _1896_ (.CLK(clk),
    .D(_0212_),
    .Q(debug_reg1[7]));
 sky130_fd_sc_hd__dfxtp_2 _1897_ (.CLK(clk),
    .D(_0213_),
    .Q(debug_reg1[8]));
 sky130_fd_sc_hd__dfxtp_2 _1898_ (.CLK(clk),
    .D(_0214_),
    .Q(debug_reg1[9]));
 sky130_fd_sc_hd__dfxtp_2 _1899_ (.CLK(clk),
    .D(_0215_),
    .Q(debug_reg1[10]));
 sky130_fd_sc_hd__dfxtp_2 _1900_ (.CLK(clk),
    .D(_0216_),
    .Q(debug_reg1[11]));
 sky130_fd_sc_hd__dfxtp_2 _1901_ (.CLK(clk),
    .D(_0217_),
    .Q(debug_reg1[12]));
 sky130_fd_sc_hd__dfxtp_2 _1902_ (.CLK(clk),
    .D(_0218_),
    .Q(debug_reg1[13]));
 sky130_fd_sc_hd__dfxtp_2 _1903_ (.CLK(clk),
    .D(_0219_),
    .Q(debug_reg1[14]));
 sky130_fd_sc_hd__dfxtp_2 _1904_ (.CLK(clk),
    .D(_0220_),
    .Q(debug_reg1[15]));
 sky130_fd_sc_hd__dfxtp_2 _1905_ (.CLK(clk),
    .D(_0221_),
    .Q(debug_reg1[16]));
 sky130_fd_sc_hd__dfxtp_2 _1906_ (.CLK(clk),
    .D(_0222_),
    .Q(debug_reg1[17]));
 sky130_fd_sc_hd__dfxtp_2 _1907_ (.CLK(clk),
    .D(_0223_),
    .Q(debug_reg1[18]));
 sky130_fd_sc_hd__dfxtp_2 _1908_ (.CLK(clk),
    .D(_0224_),
    .Q(debug_reg1[19]));
 sky130_fd_sc_hd__dfxtp_2 _1909_ (.CLK(clk),
    .D(_0225_),
    .Q(debug_reg1[20]));
 sky130_fd_sc_hd__dfxtp_2 _1910_ (.CLK(clk),
    .D(_0226_),
    .Q(debug_reg1[21]));
 sky130_fd_sc_hd__dfxtp_2 _1911_ (.CLK(clk),
    .D(_0227_),
    .Q(debug_reg1[22]));
 sky130_fd_sc_hd__dfxtp_2 _1912_ (.CLK(clk),
    .D(_0228_),
    .Q(debug_reg1[23]));
 sky130_fd_sc_hd__dfxtp_2 _1913_ (.CLK(clk),
    .D(_0229_),
    .Q(debug_reg1[24]));
 sky130_fd_sc_hd__dfxtp_2 _1914_ (.CLK(clk),
    .D(_0230_),
    .Q(debug_reg1[25]));
 sky130_fd_sc_hd__dfxtp_2 _1915_ (.CLK(clk),
    .D(_0231_),
    .Q(debug_reg1[26]));
 sky130_fd_sc_hd__dfxtp_2 _1916_ (.CLK(clk),
    .D(_0232_),
    .Q(debug_reg1[27]));
 sky130_fd_sc_hd__dfxtp_2 _1917_ (.CLK(clk),
    .D(_0233_),
    .Q(debug_reg1[28]));
 sky130_fd_sc_hd__dfxtp_2 _1918_ (.CLK(clk),
    .D(_0234_),
    .Q(debug_reg1[29]));
 sky130_fd_sc_hd__dfxtp_2 _1919_ (.CLK(clk),
    .D(_0235_),
    .Q(debug_reg1[30]));
 sky130_fd_sc_hd__dfxtp_2 _1920_ (.CLK(clk),
    .D(_0236_),
    .Q(debug_reg1[31]));
 sky130_fd_sc_hd__dfxtp_2 _1921_ (.CLK(clk),
    .D(_0237_),
    .Q(\forwarding_unit.reg_write_mem ));
 sky130_fd_sc_hd__dfxtp_2 _1922_ (.CLK(clk),
    .D(_0238_),
    .Q(id_reg_write));
 sky130_fd_sc_hd__dfxtp_2 _1923_ (.CLK(clk),
    .D(_0239_),
    .Q(\id_alu_src[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1924_ (.CLK(clk),
    .D(_0240_),
    .Q(\id_ex_rs1_data[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1925_ (.CLK(clk),
    .D(_0241_),
    .Q(\id_ex_rs1_data[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1926_ (.CLK(clk),
    .D(_0242_),
    .Q(\id_ex_rs1_data[2] ));
 sky130_fd_sc_hd__dfxtp_2 _1927_ (.CLK(clk),
    .D(_0243_),
    .Q(\id_ex_rs1_data[3] ));
 sky130_fd_sc_hd__dfxtp_2 _1928_ (.CLK(clk),
    .D(_0244_),
    .Q(\id_ex_rs1_data[4] ));
 sky130_fd_sc_hd__dfxtp_2 _1929_ (.CLK(clk),
    .D(_0245_),
    .Q(\id_ex_rs1_data[5] ));
 sky130_fd_sc_hd__dfxtp_2 _1930_ (.CLK(clk),
    .D(_0246_),
    .Q(\id_ex_rs1_data[6] ));
 sky130_fd_sc_hd__dfxtp_2 _1931_ (.CLK(clk),
    .D(_0247_),
    .Q(\id_ex_rs1_data[7] ));
 sky130_fd_sc_hd__dfxtp_2 _1932_ (.CLK(clk),
    .D(_0248_),
    .Q(\id_ex_rs1_data[8] ));
 sky130_fd_sc_hd__dfxtp_2 _1933_ (.CLK(clk),
    .D(_0249_),
    .Q(\id_ex_rs1_data[9] ));
 sky130_fd_sc_hd__dfxtp_2 _1934_ (.CLK(clk),
    .D(_0250_),
    .Q(\id_ex_rs1_data[10] ));
 sky130_fd_sc_hd__dfxtp_2 _1935_ (.CLK(clk),
    .D(_0251_),
    .Q(\id_ex_rs1_data[11] ));
 sky130_fd_sc_hd__dfxtp_2 _1936_ (.CLK(clk),
    .D(_0252_),
    .Q(\id_ex_rs1_data[12] ));
 sky130_fd_sc_hd__dfxtp_2 _1937_ (.CLK(clk),
    .D(_0253_),
    .Q(\id_ex_rs1_data[13] ));
 sky130_fd_sc_hd__dfxtp_2 _1938_ (.CLK(clk),
    .D(_0254_),
    .Q(\id_ex_rs1_data[14] ));
 sky130_fd_sc_hd__dfxtp_2 _1939_ (.CLK(clk),
    .D(_0255_),
    .Q(\id_ex_rs1_data[15] ));
 sky130_fd_sc_hd__dfxtp_2 _1940_ (.CLK(clk),
    .D(_0256_),
    .Q(\id_ex_rs1_data[16] ));
 sky130_fd_sc_hd__dfxtp_2 _1941_ (.CLK(clk),
    .D(_0257_),
    .Q(\id_ex_rs1_data[17] ));
 sky130_fd_sc_hd__dfxtp_2 _1942_ (.CLK(clk),
    .D(_0258_),
    .Q(\id_ex_rs1_data[18] ));
 sky130_fd_sc_hd__dfxtp_2 _1943_ (.CLK(clk),
    .D(_0259_),
    .Q(\id_ex_rs1_data[19] ));
 sky130_fd_sc_hd__dfxtp_2 _1944_ (.CLK(clk),
    .D(_0260_),
    .Q(\id_ex_rs1_data[20] ));
 sky130_fd_sc_hd__dfxtp_2 _1945_ (.CLK(clk),
    .D(_0261_),
    .Q(\id_ex_rs1_data[21] ));
 sky130_fd_sc_hd__dfxtp_2 _1946_ (.CLK(clk),
    .D(_0262_),
    .Q(\id_ex_rs1_data[22] ));
 sky130_fd_sc_hd__dfxtp_2 _1947_ (.CLK(clk),
    .D(_0263_),
    .Q(\id_ex_rs1_data[23] ));
 sky130_fd_sc_hd__dfxtp_2 _1948_ (.CLK(clk),
    .D(_0264_),
    .Q(\id_ex_rs1_data[24] ));
 sky130_fd_sc_hd__dfxtp_2 _1949_ (.CLK(clk),
    .D(_0265_),
    .Q(\id_ex_rs1_data[25] ));
 sky130_fd_sc_hd__dfxtp_2 _1950_ (.CLK(clk),
    .D(_0266_),
    .Q(\id_ex_rs1_data[26] ));
 sky130_fd_sc_hd__dfxtp_2 _1951_ (.CLK(clk),
    .D(_0267_),
    .Q(\id_ex_rs1_data[27] ));
 sky130_fd_sc_hd__dfxtp_2 _1952_ (.CLK(clk),
    .D(_0268_),
    .Q(\id_ex_rs1_data[28] ));
 sky130_fd_sc_hd__dfxtp_2 _1953_ (.CLK(clk),
    .D(_0269_),
    .Q(\id_ex_rs1_data[29] ));
 sky130_fd_sc_hd__dfxtp_2 _1954_ (.CLK(clk),
    .D(_0270_),
    .Q(\id_ex_rs1_data[30] ));
 sky130_fd_sc_hd__dfxtp_2 _1955_ (.CLK(clk),
    .D(_0271_),
    .Q(\id_ex_rs1_data[31] ));
 sky130_fd_sc_hd__dfxtp_2 _1956_ (.CLK(clk),
    .D(_0272_),
    .Q(\id_ex_immediate[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1957_ (.CLK(clk),
    .D(_0273_),
    .Q(\id_ex_immediate[0] ));
 sky130_fd_sc_hd__dfxtp_2 _1958_ (.CLK(clk),
    .D(_0274_),
    .Q(\id_ex_immediate[3] ));
 sky130_fd_sc_hd__dfxtp_2 _1959_ (.CLK(clk),
    .D(_0275_),
    .Q(instruction_debug[7]));
 sky130_fd_sc_hd__dfxtp_2 _1960_ (.CLK(clk),
    .D(_0276_),
    .Q(instruction_debug[15]));
 sky130_fd_sc_hd__dfxtp_2 _1961_ (.CLK(clk),
    .D(_0277_),
    .Q(instruction_debug[22]));
 sky130_fd_sc_hd__dfxtp_2 _1962_ (.CLK(clk),
    .D(_0278_),
    .Q(instruction_debug[21]));
 sky130_fd_sc_hd__conb_1 _1963_ (.HI(instruction_debug[0]));
 sky130_fd_sc_hd__conb_1 _1964_ (.HI(instruction_debug[1]));
 sky130_fd_sc_hd__conb_1 _1965_ (.HI(instruction_debug[4]));
 sky130_fd_sc_hd__conb_1 _1966_ (.LO(instruction_debug[2]));
 sky130_fd_sc_hd__conb_1 _1967_ (.LO(instruction_debug[3]));
 sky130_fd_sc_hd__conb_1 _1968_ (.LO(instruction_debug[6]));
 sky130_fd_sc_hd__conb_1 _1969_ (.LO(instruction_debug[9]));
 sky130_fd_sc_hd__conb_1 _1970_ (.LO(instruction_debug[10]));
 sky130_fd_sc_hd__conb_1 _1971_ (.LO(instruction_debug[11]));
 sky130_fd_sc_hd__conb_1 _1972_ (.LO(instruction_debug[12]));
 sky130_fd_sc_hd__conb_1 _1973_ (.LO(instruction_debug[13]));
 sky130_fd_sc_hd__conb_1 _1974_ (.LO(instruction_debug[14]));
 sky130_fd_sc_hd__conb_1 _1975_ (.LO(instruction_debug[16]));
 sky130_fd_sc_hd__conb_1 _1976_ (.LO(instruction_debug[17]));
 sky130_fd_sc_hd__conb_1 _1977_ (.LO(instruction_debug[18]));
 sky130_fd_sc_hd__conb_1 _1978_ (.LO(instruction_debug[19]));
 sky130_fd_sc_hd__conb_1 _1979_ (.LO(instruction_debug[24]));
 sky130_fd_sc_hd__conb_1 _1980_ (.LO(instruction_debug[25]));
 sky130_fd_sc_hd__conb_1 _1981_ (.LO(instruction_debug[26]));
 sky130_fd_sc_hd__conb_1 _1982_ (.LO(instruction_debug[27]));
 sky130_fd_sc_hd__conb_1 _1983_ (.LO(instruction_debug[28]));
 sky130_fd_sc_hd__conb_1 _1984_ (.LO(instruction_debug[29]));
 sky130_fd_sc_hd__conb_1 _1985_ (.LO(instruction_debug[30]));
 sky130_fd_sc_hd__conb_1 _1986_ (.LO(instruction_debug[31]));
 sky130_fd_sc_hd__conb_1 _1987_ (.LO(pc_current[0]));
 sky130_fd_sc_hd__conb_1 _1988_ (.LO(pc_current[1]));
 sky130_fd_sc_hd__buf_2 _1989_ (.A(instruction_debug[15]),
    .X(instruction_debug[5]));
 sky130_fd_sc_hd__buf_2 _1990_ (.A(instruction_debug[21]),
    .X(instruction_debug[8]));
 sky130_fd_sc_hd__buf_2 _1991_ (.A(instruction_debug[22]),
    .X(instruction_debug[20]));
 sky130_fd_sc_hd__buf_2 _1992_ (.A(mem_wb_valid),
    .X(pipeline_state[0]));
 sky130_fd_sc_hd__buf_2 _1993_ (.A(ex_mem_valid),
    .X(pipeline_state[1]));
 sky130_fd_sc_hd__buf_2 _1994_ (.A(id_ex_valid),
    .X(pipeline_state[2]));
 sky130_fd_sc_hd__buf_2 _1995_ (.A(if_id_valid),
    .X(pipeline_state[3]));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Left_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Left_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Left_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Left_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Left_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Left_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Left_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Left_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2171 ();
endmodule
